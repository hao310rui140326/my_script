module test_top(/*AUTOARG*/
   );

output   test_o ;



/*AUTOOUTPUT*/
/*AUTOINPUT*/
/*AUTOWIRE*/


/*test  AUTO_TEMPLATE( .o(o[@]),  );*/

test test0 (
/*AUTOINST*/
);


test test1 (
/*AUTOINST*/
);


test test2 (
/*AUTOINST*/
);

endmodule





