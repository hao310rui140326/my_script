 module OIIOlIO0ooOLLoll0il0IlOloL0oOIlII ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO , Oo0LLillol0loLIo0iOl0oOLlIOlILoIO , OoOi0O0oOoL0looLo0IoOllOOILiLooLl , OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI , OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII , OOLOoolOi0LIo0olO0loLllIlllIiiIiI , OOOLiLOilooIi0Iio00ilILoLIILOoOoI , OLLOooI0ILL00ILloiliILLLiioooLliI , OILoli0OIOIIOI0OiliOo0i0OLoliOOiI , O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI , O0I0oI0I000LllOOI0L0lOlIl000LIioO , OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI , OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 , OOooLlloIiioOOO0LLILl0liiillLILol , OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo , OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI , OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 , OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol , OloliIooiiLI0IIlOiL0LLlioILLllL0L , O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO , OioILlIiO0000OoolooO00loIOIloLIoI , OLOl0000OLooLIIo0lIOIOI0lILioolOl , OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII , OoIolLlOIIoIoi00lloLlIoI0lo0iILol , OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI , OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo , OOIIloOlOILliIOILOIOiIlooIOOIL0oO , OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io , OiLOo0loOI00OL0Ooio0OIIlOLiooLOII , OlLilll0ilOLI0IIoO0li0l0OlO00oLIO , O0liLooiLliIoLOllliIlo0ILo0I0oOOl , O0i00oOl00OoIIOIil0LLOi0looIOIL00 );
 parameter OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL = 5'd0 ;
 parameter Oo0oIiiLoLI0IOiI0lloIOOollollIIlL = 5'd1 ;
 parameter OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO = 5'd4 ;
 parameter OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo = 5'd5 ;
 parameter OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo = 5'd6 ;
 parameter OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 = 5'd7 ;
 parameter OllIlooiolLL00OiIIiOO0iOOiIlLLOoi = 5'd8 ;
 parameter OiilO0lI0iIIOio0IIiiOoIoioLL00oOO = 5'd22 ;
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input [15:0] OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 input OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ;
 input [ 3:0] OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 input OOLOoolOi0LIo0olO0loLllIlllIiiIiI ;
 input OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 input [63:0] OLLOooI0ILL00ILloiliILLLiioooLliI ;
 input [ 2:0] OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 input [15:0] O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ;
 input O0I0oI0I000LllOOI0L0lOlIl000LIioO ;
 output OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ;
 input OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 output OOooLlloIiioOOO0LLILl0liiillLILol ;
 output [15:0] OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ;
 output [31:0] Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 output Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ;
 output OoOi0O0oOoL0looLo0IoOllOOILiLooLl ;
 output [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 output [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 output [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 output [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 output [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 output [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 output [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 output [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 output [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 output [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 output [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 output [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 output [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 output [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 output [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 output [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 output O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 wire [31:0] Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 reg [31:0] OlOLilIOoLLlOiLloiOIl00OLLiILiiIo ;
 reg OoOi0O0oOoL0looLo0IoOllOOILiLooLl ;
 reg Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ;
 reg [ 5:0] Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ;
 reg O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ;
 wire [191:0] O0lOIlooLi0lilOllLlilIo00iOLiOLLo ;
 wire [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 wire [15:0] OILIloOoilLIL00IIOoOilLOO0L0iiIOO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:112+64];
 wire [15:0] O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 96+64];
 wire [31:0] O0oLLi0Ill00l0lioiLioiooIllloIiIl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 64+64];
 wire [15:0] Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:112+64];
 wire [31:0] OlO0Oo0looiIoIiL0liIllLLLL0o00i0L = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 80+64];
 wire [31:0] O0o0loiLIOlLoi0iOIolL0LoOILoilLLl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:96+64] ;
 wire [15:0] Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64:80+64] ;
 wire [15:0] OiO0oiLLillil0LLLOLo0OoiiOLLIILiI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 79+64:64+64] ;
 wire [15:0] OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:112+64];
 wire [15:0] OOioILiL0oiO0OIlLLOLLi0O0oOOIlIlI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 96+64];
 wire [15:0] OOiLiOlo0ioloILilO0IlILL0o0iiLiOI = 16'd81 ;
 reg [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 reg [2 :0] OOOi0LIiLLOLIoliiOlolloOli0oLLioi ;
 reg [15:0] OILLIiOoiIOiIil0OLOLLiIIllIlOLilI ;
 reg [15:0] OLIiiio00OOiooIiolIO0ooLl0OlIoloI ;
 reg [15:0] OliiLIIliIO0OIloloLiiI0ilOILLILOI ;
 reg [15:0] OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo ;
 reg [15:0] OLOlIOIOOlLOII0OLL0oiL0I0O0IilloL ;
 wire [11:0] O0oioIoloolL0oiioLILllioiO0oliIOl ;
 wire [ 3:0] Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 assign O0oioIoloolL0oiioLILllioiO0oliIOl = OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo[15:4] ;
 assign Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi = OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo[ 3:0] ;
 reg [11:0] OLIo0LL0IiLIOliLL00I0LO00IllOOllo ;
 reg [15:0] Oi0ILolLOL0li0iLIolliilIlLlloolO0 ;
 reg [15:0] OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ;
 reg OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL ;
 reg OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ;
 wire OIlii0Io00iIi0iIOilOOoollO0iI0lol = OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 reg [ 4:0] OOLIiil0IlIllLollIl0LIilliOI0iolo ;
 reg [ 4:0] OL0II0lIOioLIIOLlLILoioOiOLLlLLLL ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLIiil0IlIllLollIl0LIilliOI0iolo <= 5'd0 ;
 end
 else if (OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI||OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OOLIiil0IlIllLollIl0LIilliOI0iolo <= 5'd0 ;
 end
 else begin
 OOLIiil0IlIllLollIl0LIilliOI0iolo <= OL0II0lIOioLIIOLlLILoioOiOLLlLLLL ;
 end
 end
 wire Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL );
 wire Olo0LI0lIlil0IIloOOIoi0L0LOoIIoOl = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== Oo0oIiiLoLI0IOiI0lloIOOollollIIlL );
 wire O0LO0iloLil0LI0IOiOolIoioLOOIOLiO = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO );
 wire OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo );
 wire OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo );
 wire OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 );
 wire OOIIIOLL0O000ioLliOIoOii0LiI0lOoo = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OllIlooiolLL00OiIIiOO0iOOiIlLLOoi );
 always@ ( * ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OOLIiil0IlIllLollIl0LIilliOI0iolo;
 case(OOLIiil0IlIllLollIl0LIilliOI0iolo) OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL : begin
 if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = Oo0oIiiLoLI0IOiI0lloIOOollollIIlL ;
 end
 end
 Oo0oIiiLoLI0IOiI0lloIOOollollIIlL : begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) begin
 if ((OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiilO0lI0iIIOio0IIiiOoIoioLL00oOO ;
 end
 end
 end
 OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO : begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd6 ) begin
 if ( ( Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) &&(OlO0Oo0looiIoIiL0liIllLLLL0o00i0L==32'h0000_5902) ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiilO0lI0iIIOio0IIiiOoIoioLL00oOO ;
 end
 end
 end
 OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) begin
 if (Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI<=16'h0001) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo ;
 end
 end
 end
 /* OoIlLOiLLl0Il0Ili0Lo0ooLloO00oILL : begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi>=(OlI0LilLLoO0OiiLioLoIIILooLIlILOi-1'b1)) ) begin
 if ( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0==4'd0 ) begin
 if ( OolIOLOooiLLIllI0LOLIolllLoilolIl<(16'd16+ OOiLiOlo0ioloILilO0IlILL0o0iiLiOI ) ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = FIR_R_DSYNC_STATE ;
 end
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = O0IloLIOl0I0oli0IOIoOO0lOolioolIl ;
 end
 end
 end
 O0IloLIOl0I0oli0IOIoOO0lOolioolIl: begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ) begin
 if ( OolIOLOooiLLIllI0LOLIolllLoilolIl<( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 + OOiLiOlo0ioloILilO0IlILL0o0iiLiOI )) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = FIR_R_DSYNC_STATE ;
 end
 end
 end
 */ OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4 )begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 ;
 end
 end
 OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 : begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) )begin
 if (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo ;
 end
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OllIlooiolLL00OiIIiOO0iOOiIlLLOoi ;
 end
 end
 end
 OllIlooiolLL00OiIIiOO0iOOiIlLLOoi : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo ;
 end
 end
 end
 /* OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L : begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl==16'd0) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else if (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ? O0Il0i0oII0Lil0IooLoIIliOoOI0oiO0 : FIR_RSC_SEGMT_H_STATE ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiIoi0liOllioIL0IilOLIOIOIiILiioI ;
 end
 end
 */ /* O0Il0i0oII0Lil0IooLoIIliOoOI0oiO0 : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 FIR_RSC_SEGMT_H_STATE : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 */ /* FIR_RSC_SEGMT_STATE : begin
 if ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)&&(OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd16)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = FIR_RSC_SEGMT_END_STATE ;
 end
 end
 FIR_RSC_SEGMT_END_STATE : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 O0OiiIi0olIo0IIL0O0OIIolIiIOLllO0 : begin
 if ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)&&(OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd16)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OILlioiLloo0oIiI0o0ILOIIiO0IoiOil ;
 end
 end
 OILlioiLloo0oIiI0o0ILOIIiO0IoiOil : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 */ OiilO0lI0iIIOio0IIiiOoIoioLL00oOO : begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 default : begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 endcase end
 /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 <= 1'd0 ;
 sc_frame_flag <= 1'd0 ;
 end
 else if ( O0LO0iloLil0LI0IOiOolIoioLOOIOLiO ) begin
 OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 <= (Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==16'h03e9) ;
 sc_frame_flag <= (Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==16'h1389) ;
 end
 end
 */ /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0IIOiLIOiIi0Ol0000ilIill0II0OilI <= 16'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI&&~tcp_scmatch_flag) begin
 O0IIOiLIOiIi0Ol0000ilIill0II0OilI <= OilOOioILlOIIOL0iioIOIi0oloooOoLl - 16'd22 ;
 end
 else if ( fir_r_dsync_st || OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) begin
 O0IIOiLIOiIi0Ol0000ilIill0II0OilI <= O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo - 16'd22 ;
 end
 end
 */ /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= 16'd0 ;
 end
 else if ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= (OIIOLLOIlOlLoi0oiOioLilOiioiiliLO - O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI - OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII - 16'd8) ;
 end
 else if ( ( fir_r_dsync_st || OlliILlLOilOl0LO0O0OilooiIIiOi0Ll) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if (O0LO0iloLil0LI0IOiOolIoioLOOIOLiO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd6) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd6 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd12) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd12 ;
 end
 else if (OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd4) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd4 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd16 ;
 end
 else if (OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 end
 else if ( (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl || fir_r_sccut_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if ( (OIoIooIolOilIOlooOlOIIOoilLioOIIO || fir_r_sccut_end_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ( (O0oill0llILOilo0i0LIoOLIoolL0Il0o || fir_r_sccuth_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ((OiL0LolLLIOlliloII00llOil0oIlOiIo) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if ((O0llIOIliLOO0iiOoO0OO0lIOloLoII0I) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 end
 else if ((fir_r_scrcut_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if ((fir_r_scrcut_end_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=sub_sccut_len_reg) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - sub_sccut_len_reg ;
 end
 end
 */ reg [3:0] OLliloOlllioIloi0iiloI00oOLoOoO0L ;
 reg [3:0] Oi0llIo0lIioooLLII00oOiO0LI0LILio ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd0 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= 4'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd0 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= 4'd0 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO&&( OOLIiil0IlIllLollIl0LIilliOI0iolo>= OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ) ) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd0 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= 4'd0 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO&&( OOLIiil0IlIllLollIl0LIilliOI0iolo== OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ) ) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd0 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= 4'd0 ;
 end
 else if (OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL&& ( OOLIiil0IlIllLollIl0LIilliOI0iolo>= OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ) ) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd0 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= 4'd0 ;
 end
 else if (OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL && (OLliloOlllioIloi0iiloI00oOLoOoO0L>=4'd7) ) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd0 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= 4'd0 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO ) begin
 OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL <= 1'd1 ;
 OLliloOlllioIloi0iiloI00oOLoOoO0L <= OLliloOlllioIloi0iiloI00oOLoOoO0L + 4'd1 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oi0llIo0lIioooLLII00oOiO0LI0LILio <= 1'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 Oi0llIo0lIioooLLII00oOiO0LI0LILio <= 1'd0 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO ) begin
 Oi0llIo0lIioooLLII00oOiO0LI0LILio <= Oi0llIo0lIioooLLII00oOiO0LI0LILio + 1'd1 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd1 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO&&( OOLIiil0IlIllLollIl0LIilliOI0iolo>= OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ) ) begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd1 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO&&( OOLIiil0IlIllLollIl0LIilliOI0iolo== OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ) ) begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd1 ;
 end
 else if (OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL&& ( OOLIiil0IlIllLollIl0LIilliOI0iolo>= OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ) ) begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd1 ;
 end
 else if (OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL && (OLliloOlllioIloi0iiloI00oOLoOoO0L>=4'd7) ) begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd1 ;
 end
 else begin
 OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOOi0LIiLLOLIoliiOlolloOli0oLLioi <= 3'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li ) begin
 OOOi0LIiLLOLIoliiOlolloOli0oLLioi <= (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) ? OOOi0LIiLLOLIoliiOlolloOli0oLLioi + 1'd1 : OOOi0LIiLLOLIoliiOlolloOli0oLLioi ;
 end
 else begin
 OOOi0LIiLLOLIoliiOlolloOli0oLLioi <= 3'd0 ;
 end
 end
 reg OIoOolllLOOiliOLL0oOLo0LLloIOOi0l ;
 reg OOoIliOliILLi0IiIlILLo00iLoLiloIl ;
 reg OIIILoOLllIiLloiiIoiiLooiiI00Oii0 ;
 reg OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 ;
 reg OI00liOIoliolOollOLoioOLooloiloI0 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo <= 16'd0 ;
 OLOlIOIOOlLOII0OLL0oiL0I0O0IilloL <= 16'd0 ;
 OIoOolllLOOiliOLL0oOLo0LLloIOOi0l <= 1'd0 ;
 OOoIliOliILLi0IiIlILLo00iLoLiloIl <= 1'd0 ;
 OIIILoOLllIiLloiiIoiiLooiiI00Oii0 <= 1'd0 ;
 end
 else if ( OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4) ) begin
 OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo <= OOioILiL0oiO0OIlLLOLLi0O0oOOIlIlI ;
 OLOlIOIOOlLOII0OLL0oiL0I0O0IilloL <= OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL ;
 OIoOolllLOOiliOLL0oOLo0LLloIOOi0l <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2439) ;
 OOoIliOliILLi0IiIlILLo00iLoLiloIl <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2433) ;
 OIIILoOLllIiLloiiIoiiLooiiI00Oii0 <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2434) ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 <= 1'd0 ;
 OI00liOIoliolOollOLoioOLooloiloI0 <= 1'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 <= 1'd0 ;
 OI00liOIoliolOollOLoioOLooloiloI0 <= 1'd0 ;
 end
 else if ( OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4) ) begin
 OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2433) ? 1'd1 : OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 ;
 OI00liOIoliolOollOLoioOLooloiloI0 <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2434) ? 1'd1 : OI00liOIoliolOollOLoioOLooloiloI0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OILLIiOoiIOiIil0OLOLLiIIllIlOLilI <= 16'd0 ;
 OLIiiio00OOiooIiolIO0ooLl0OlIoloI <= 16'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) ) begin
 OILLIiOoiIOiIil0OLOLLiIIllIlOLilI <= Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI ;
 OLIiiio00OOiooIiolIO0ooLl0OlIoloI <= OiO0oiLLillil0LLLOLo0OoiiOLLIILiI ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OliiLIIliIO0OIloloLiiI0ilOILLILOI <= 16'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OliiLIIliIO0OIloloLiiI0ilOILLILOI <= 16'd0 ;
 end
 else if ( OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4 ) ) begin
 OliiLIIliIO0OIloloLiiI0ilOILLILOI <= OliiLIIliIO0OIloloLiiI0ilOILLILOI + 1'd1 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 /* else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI&&~tcp_scmatch_flag && OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd6 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OI00OiLolooiIIiiILoIliO0O0loolIlI && OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 */ else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OIlii0Io00iIi0iIOilOOoollO0iI0lol && (OILoli0OIOIIOI0OiliOo0i0OLoliOOiI==3'd0) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 /* else if (OiL0LolLLIOlliloII00llOil0oIlOiIo) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l<=16'd16) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]))) ? Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] - 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]))) ? 1'd1 : 1'd0;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I && ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8))) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8))) ? 1'd1 : 1'd0 ;
 end
 else if (fir_r_scrcut_st) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (sub_sccut_len_reg<=16'd16) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(sub_sccut_len_reg[5:0]))) ? sub_sccut_len_reg[5:0] - 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(sub_sccut_len_reg[5:0]))) ? 1'd1 : 1'd0;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (fir_r_scrcut_end_st && ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=sub_sccut_len_reg[5:0] ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(sub_sccut_len_reg[5:0]+6'd8))) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(sub_sccut_len_reg[5:0]+6'd8))) ? 1'd1 : 1'd0 ;
 end
 */ else if (Olo0LI0lIlil0IIloOOIoi0L0LOoIIoOl ) begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd14)|| (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd6)) ? 6'd6 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd14)|| (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd6)) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol && ((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd8) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 /* else if (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) begin
 if ( (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && (OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0||sc_frame_flag) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 if ((OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd4 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 */ else if (O0LO0iloLil0LI0IOiOolIoioLOOIOLiO) begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd6 ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd18)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd2-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd12))) ? 6'd12 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd18)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd2-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd12))) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd6)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd6 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol-6'd4-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd4))) ? 6'd4 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&((O0IOooLliOlIllOliILoolIIoIiO0Ilol-6'd4-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd4))) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd12) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd12 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 /* else if ( Oo0LiLOLOIi0lLoOlLLiIoo00lLlloOlO ) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi>=(OlI0LilLLoO0OiiLioLoIIILooLIlILOi-1'b1)) ) begin
 if ( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0==4'd0 ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd24)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16))) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd24)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16))) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd16+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0)))) ? Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd16+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0)))) ? 1'd1 : 1'd0 ;
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd16 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OLIoo0OL0oo0iloLooi0iIIoLLOlIILIL) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0)))) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0)))) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 */ else if (OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4 )begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd4-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd16) )) ? 6'd16 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd4-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd16) )) ? 1'd1 : 1'd0 ;
 end
 else if ( OIlii0Io00iIi0iIOilOOoollO0iI0lol && ((O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd4) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd4 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) )begin
 if (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI<OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)|| (OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ((O0IOooLliOlIllOliILoolIIoIiO0Ilol-6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd4) ) ) ? 6'd4 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)|| (OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ((O0IOooLliOlIllOliILoolIIoIiO0Ilol-6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>=6'd4) ) ) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd16+Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol && ((O0IOooLliOlIllOliILoolIIoIiO0Ilol-6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)>= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+OILoli0OIOIIOI0OiliOo0i0OLoliOOiI)) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? 6'd0 : 6'd16 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? 1'd0 : 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo ) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 else begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd4+Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd4 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if ( OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(OILoli0OIOIIOI0OiliOo0i0OLoliOOiI<=6'd4 ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd4 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if ( OIlii0Io00iIi0iIOilOOoollO0iI0lol && ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol + 6'd8) >= (6'd4 + OILoli0OIOIIOI0OiliOo0i0OLoliOOiI + Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi )) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd4 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8-OILoli0OIOIIOI0OiliOo0i0OLoliOOiI) >= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 /* else if (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl==16'd0) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 else if (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= OolIOLOooiLLIllI0LOLIolllLoilolIl[5:0] ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 end
 */ /* else if (fir_r_sccut_st || OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) begin
 if ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)&&(OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd16)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(OolIOLOooiLLIllI0LOLIolllLoilolIl))||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? (OolIOLOooiLLIllI0LOLIolllLoilolIl[5:0]-6'd8) : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(OolIOLOooiLLIllI0LOLIolllLoilolIl))||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 */ else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 wire [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 wire [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 reg [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 wire [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 wire [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 reg [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 reg [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 reg [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 reg [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 reg [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 reg [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 reg [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 reg [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 reg [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 reg [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 reg [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 reg O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol <= 32'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) ) begin
 OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol <= {O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[7:0],O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[15:8],O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[23:16],O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[31:24]} ;
 end
 end
 wire [127: 0] OILiOOlOoOl0OiO0OlOoOliIILlliioOl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 64] ;
 wire [ 47: 0] OIIooioLOLO0OIiOiiiooOOIOI0OollII = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:80+64] ;
 wire [ 71: 0] OIlIOllOoilOIlI0OLLoL0l00l0ilooIi = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 79+64: 8+64] ;
 wire [ 7: 0] OiLOLi0io00oIo00Io0lLlLIL0lioiI00 = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 7+64: 64] ;
 wire [ 63: 0] OOILIooliL0iOIOlilO0OiLlLoLIiLOil = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:64+64] ;
 wire [ 31: 0] OOIliIiiiilolLLLLLoi0IlLoilIIOiII = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64:32+64] ;
 wire [ 63: 0] Oo0OioiiiiIiloIIL0ILILoliiO0iooOL = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 64+64] ;
 wire [ 31: 0] OiILllOLOIIl00ooOllolL0OiIIIIOlL0 = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64: 32+64] ;
 wire [ 31: 0] OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 31+64: 64] ;
 wire [ 31: 0] OlooLooOLllollooO0LLIIOilii0o0OlO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 96+64] ;
 wire [ 63: 0] Ol0oii0iIi0Ioo0loOil0000LooOL0OOl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 32+64] ;
 wire [ 63: 0] OOIOIOIOooiooiilLoOIoL0olL0O0o0Il = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 64+64] ;
 wire [ 31: 0] O0OLLl000lO0LIi0o00iolO0ILoIlOi0O = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64: 32+64] ;
 wire [ 31: 0] OilOOoIIOl0liLOilL0o0LiliIioOLOiI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 31+64: 64] ;
 wire [ 31: 0] OolOIilLOLOLLLiIoOlloool0lolooiO0 = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 96+64] ;
 wire [ 31: 0] OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 64+64] ;
 assign OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI = {8'h53,8'h51,8'h00} ;
 assign OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 = 8'h31 ;
 assign OloliIooiiLI0IIlOiL0LLlioILLllL0L = 8'h30 ;
 assign O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO = 32'd0 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OioILlIiO0000OoolooO00loIOIloLIoI <= 176'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OioILlIiO0000OoolooO00loIOIloLIoI <= 176'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OioILlIiO0000OoolooO00loIOIloLIoI[175:48] <= OILiOOlOoOl0OiO0OlOoOliIILlliioOl ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd1) ) begin
 OioILlIiO0000OoolooO00loIOIloLIoI[47: 0] <= OIIooioLOLO0OIiOiiiooOOIOI0OollII ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl <= 72'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl <= 72'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd1) ) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl[71:64] <= OiLOLi0io00oIo00Io0lLlLIL0lioiI00 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd2) ) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl[63: 0] <= OOILIooliL0iOIOlilO0OiLlLoLIiLOil ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd2) ) begin
 OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII[31: 0] <= {OOIliIiiiilolLLLLLoi0IlLoilIIOiII[7:0],OOIliIiiiilolLLLLLoi0IlLoilIIOiII[15:8],OOIliIiiiilolLLLLLoi0IlLoilIIOiII[23:16],OOIliIiiiilolLLLLLoi0IlLoilIIOiII[31:24]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OoIolLlOIIoIoi00lloLlIoI0lo0iILol <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OoIolLlOIIoIoi00lloLlIoI0lo0iILol[63:0]) ) begin
 OoIolLlOIIoIoi00lloLlIoI0lo0iILol <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OoIolLlOIIoIoi00lloLlIoI0lo0iILol[63: 0] <= {Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[7:0],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[15:8],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[23:16],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[31:24],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[39:32],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[47:40],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[55:48],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[63:56]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI[31: 0] <= { OiILllOLOIIl00ooOllolL0OiIIIIOlL0[7:0],OiILllOLOIIl00ooOllolL0OiIIIIOlL0[15:8],OiILllOLOIIl00ooOllolL0OiIIIIOlL0[23:16],OiILllOLOIIl00ooOllolL0OiIIIIOlL0[31:24] } ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[63:0]) ) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[31: 0] <= { OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[7:0],OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[15:8],OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[23:16],OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[31:24] } ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) ) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[63: 32] <= { OlooLooOLllollooO0LLIIOilii0o0OlO[7:0],OlooLooOLllollooO0LLIIOilii0o0OlO[15:8],OlooLooOLllollooO0LLIIOilii0o0OlO[23:16],OlooLooOLllollooO0LLIIOilii0o0OlO[31:24] } ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOIIloOlOILliIOILOIOiIlooIOOIL0oO <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OOIIloOlOILliIOILOIOiIlooIOOIL0oO[63:0]) ) begin
 OOIIloOlOILliIOILOIOiIlooIOOIL0oO <= 'd0 ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) ) begin
 OOIIloOlOILliIOILOIOiIlooIOOIL0oO[63: 0] <= {Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[7:0],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[15:8],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[23:16],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[31:24],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[39:32],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[47:40],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[55:48],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[63:56]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io[63:0]) ) begin
 OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io[63: 0] <= {OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[7:0],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[15:8],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[23:16],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[31:24],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[39:32],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[47:40],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[55:48],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[63:56]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiLOo0loOI00OL0Ooio0OIIlOLiooLOII <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OiLOo0loOI00OL0Ooio0OIIlOLiooLOII <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OiLOo0loOI00OL0Ooio0OIIlOLiooLOII[31: 0] <= {O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[7:0],O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[15:8],O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[23:16],O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[31:24]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO ) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==3'd0) ) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[31: 0] <= {OilOOoIIOl0liLOilL0o0LiliIioOLOiI[7:0],OilOOoIIOl0liLOilL0o0LiliIioOLOiI[15:8],OilOOoIIOl0liLOilL0o0LiliIioOLOiI[23:16],OilOOoIIOl0liLOilL0o0LiliIioOLOiI[31:24] } ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) ) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[63: 0] <= ((&OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[31: 0])&&(&OolOIilLOLOLLLiIoOlloool0lolooiO0[31:0])) ? 64'd0 : { {OolOIilLOLOLLLiIoOlloool0lolooiO0[7:0],OolOIilLOLOLLLiIoOlloool0lolooiO0[15:8],OolOIilLOLOLLLiIoOlloool0lolooiO0[23:16],OolOIilLOLOLLLiIoOlloool0lolooiO0[31:24] } , OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[31:0] } ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0liLooiLliIoLOllliIlo0ILo0I0oOOl <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 O0liLooiLliIoLOllliIlo0ILo0I0oOOl <= 'd0 ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) ) begin
 O0liLooiLliIoLOllliIlo0ILo0I0oOOl[31: 0] <= {OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[7:0],OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[15:8],OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[23:16],OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[31:24]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlOLilIOoLLlOiLloiOIl00OLLiILiiIo <= 32'd0 ;
 OoOi0O0oOoL0looLo0IoOllOOILiLooLl <= 1'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi||O0LO0iloLil0LI0IOiOolIoioLOOIOLiO) begin
 OlOLilIOoLLlOiLloiOIl00OLLiILiiIo <= 32'd0 ;
 OoOi0O0oOoL0looLo0IoOllOOILiLooLl <= 1'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ) begin
 OlOLilIOoLLlOiLloiOIl00OLLiILiiIo <= O0o0loiLIOlLoi0iOIolL0LoOILoilLLl ;
 OoOi0O0oOoL0looLo0IoOllOOILiLooLl <= 1'd1 ;
 end
 else begin
 OoOi0O0oOoL0looLo0IoOllOOILiLooLl <= 1'd0 ;
 end
 end
 assign Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO = OlOLilIOoLLlOiLloiOIl00OLLiILiiIo ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li ) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) )begin
 if (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 end
 else begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 end
 else begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 end
 else begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 end
 else if (OOIIIOLL0O000ioLliOIoOii0LiI0lOoo) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 end
 else begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 end
 else begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 end
 else begin
 Oo0LLillol0loLIo0iOl0oOLlIOlILoIO <= 1'd0 ;
 end
 end
 /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo <= 32'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) ) begin
 if ( (O0o0loiLIOlLoi0iOIolL0LoOILoilLLl>OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&&OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && (Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI>16'h0001) ) begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo = O0o0loiLIOlLoi0iOIolL0LoOILoilLLl ;
 end
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 current_scid_reg <= 32'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) ) begin
 if ( (O0o0loiLIOlLoi0iOIolL0LoOILoilLLl>current_scid_reg)&&sc_frame_flag && (Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI>16'h0001) ) begin
 current_scid_reg = O0o0loiLIOlLoi0iOIolL0LoOILoilLLl ;
 end
 end
 end
 */ /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 sc_cut_flag <= 1'd0 ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) ) begin
 sc_cut_flag <= sc_frame_flag ;
 end
 else if (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL) begin
 sc_cut_flag <= sc_frame_flag && (|OolIOLOooiLLIllI0LOLIolllLoilolIl) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8) ;
 end
 else begin
 sc_cut_flag <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O <= 1'd0 ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) ) begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O <= OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 end
 else if (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL) begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O <= OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && (|OolIOLOooiLLIllI0LOLIolllLoilolIl) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8 ) ;
 end
 else begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O <= 1'd0 ;
 end
 end
 */ always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= 1'd0 ;
 end
 else if (O0I0oI0I000LllOOI0L0lOlIl000LIioO || OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI || OL0OI0o0lILOoIoIiiLiOOLIoiilo0liL ) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= 1'd0 ;
 end
 else if (OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) && (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) && (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) ) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= (OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 || OI00liOIoliolOollOLoioOLooloiloI0) ;
 end
 else if (OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) && (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) ) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= (OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 || OI00liOIoliolOollOLoioOLooloiloI0) ;
 end
 else begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= 1'd0 ;
 end
 end
 /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OL0O0IIio0loL0L0Il0li0i00lliIoOOI <= 1'd1 ;
 end
 else if (OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1)) && (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) && (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) ) begin
 OL0O0IIio0loL0L0Il0li0i00lliIoOOI <= 1'd0 ;
 end
 else if (OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) && (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) ) begin
 OL0O0IIio0loL0L0Il0li0i00lliIoOOI <= 1'd0 ;
 end
 else if ( OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL ) begin
 OL0O0IIio0loL0L0Il0li0i00lliIoOOI <= 1'd1 ;
 end
 else begin
 OL0O0IIio0loL0L0Il0li0i00lliIoOOI <= 1'd1 ;
 end
 end
 */ always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= 16'd81 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= 16'd81 ;
 end
 else if ( Olo0LI0lIlil0IIloOOIoi0L0LOoIIoOl && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo + 16'd4 ;
 end
 end
 /* always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= 16'd0 ;
 end
 else if ( O0oill0llILOilo0i0LIoOLIoolL0Il0o ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= 16'd8 ;
 end
 else if ( (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (OolIOLOooiLLIllI0LOLIolllLoilolIl>16'd8) ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo + 16'd8 ;
 end
 else if ( (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8) ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if (OiL0LolLLIOlliloII00llOil0oIlOiIo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) && (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l>16'd8) ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo + 16'd8 ;
 end
 else if (OiL0LolLLIOlliloII00llOil0oIlOiIo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l) && (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l<=16'd8) ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo + Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 st_rc_cut_cnt <= 16'd0 ;
 end
 else if ( fir_r_sccuth_st ) begin
 st_rc_cut_cnt <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && sc_frame_flag ) begin
 st_rc_cut_cnt <= 16'd8 ;
 end
 else if ( ( fir_r_sccut_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (OolIOLOooiLLIllI0LOLIolllLoilolIl>16'd8) ) begin
 st_rc_cut_cnt <= st_rc_cut_cnt + 16'd8 ;
 end
 else if ( ( fir_r_sccut_st) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8) ) begin
 st_rc_cut_cnt <= st_rc_cut_cnt + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if (fir_r_scrcut_st && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) && (sub_sccut_len_reg>16'd8) ) begin
 st_rc_cut_cnt <= st_rc_cut_cnt + 16'd8 ;
 end
 else if (fir_r_scrcut_st && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=sub_sccut_len_reg) && (sub_sccut_len_reg<=16'd8) ) begin
 st_rc_cut_cnt <= st_rc_cut_cnt + sub_sccut_len_reg ;
 end
 end
 */ /* OoLiL0iillLiLlLlO0loIIoLl0l0l0LoI sq_fir_cut_out ( .OilOIloOO0LiLoIL0IIILoIi0Loilll0I (OilOIloOO0LiLoIL0IIILoIi0Loilll0I ), .Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 (Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ), .OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O (OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ), .OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO (OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ), .OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 (OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ), .O0oill0llILOilo0i0LIoOLIoolL0Il0o (O0oill0llILOilo0i0LIoOLIoolL0Il0o ), .OlliILlLOilOl0LO0O0OilooiIIiOi0Ll (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ), .OOLoL0looIOoioIoOooIoLIiIiLiLoiOl (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ), .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ), .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl ), .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 (OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ), .O0lOIlooLi0lilOllLlilIo00iOLiOLLo (O0lOIlooLi0lilOllLlilIo00iOLiOLLo ), .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo ), .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) );
 OoLiL0iillLiLlLlO0loIIoLl0l0l0LoI sc_fir_cut_out ( .OilOIloOO0LiLoIL0IIILoIi0Loilll0I (sc_rx_start ), .Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 (sc_rx_end ), .OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O (sc_rx_valid ), .OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO (sc_rx_data ), .OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 (sc_rx_empty ), .O0oill0llILOilo0i0LIoOLIoolL0Il0o (fir_r_sccuth_st ), .OlliILlLOilOl0LO0O0OilooiIIiOi0Ll (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ), .OOLoL0looIOoioIoOooIoLIiIiLiLoiOl (fir_r_sccut_st ), .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ), .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl ), .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 (sc_frame_flag ), .O0lOIlooLi0lilOllLlilIo00iOLiOLLo (O0lOIlooLi0lilOllLlilIo00iOLiOLLo ), .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo ), .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) );
 */ OLiIILolLli0LiLoOOo0lIlOiOoO0lioL OLiIILolLli0LiLoOOo0lIlOiOoO0lioL ( .OOLIiil0IlIllLollIl0LIilliOI0iolo (OOLIiil0IlIllLollIl0LIilliOI0iolo ) , .O0il0IO0olIoLiOIL0000lo0OoliIL0Ll (OOooLlloIiioOOO0LLILl0liiillLILol ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII (4'd0 ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI (OOLOoolOi0LIo0olO0loLllIlllIiiIiI ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI (OOOLiLOilooIi0Iio00ilILoLIILOoOoI ) , .OLLOooI0ILL00ILloiliILLLiioooLliI (OLLOooI0ILL00ILloiliILLLiioooLliI ) , .OL0O0IIio0loL0L0Il0li0i00lliIoOOI (1'd1 ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI (OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ) , .Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ) , .O0lOIlooLi0lilOllLlilIo00iOLiOLLo (O0lOIlooLi0lilOllLlilIo00iOLiOLLo ) , .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ) , .Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl (Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ) , .O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI (O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ) , .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) );
 endmodule
 module OiI00lI0lL0IoLLLlLoioLlOIOOiOiiIi ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L , OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl , OoIolioOL0iLLOLloI00iIILLiiL0Ooil , Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 , OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI , OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 , OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI , OilOOo00lLiOOoiO0ii0oo0oOliOollii , OolIOLOooiLLIllI0LOLIolllLoilolIl , O0IOooLliOlIllOliILoolIIoIiO0Ilol , O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo , OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 , OILIloOoilLIL00IIOoOilLOO0L0iiIOO , O0oLLi0Ill00l0lioiLioiooIllloIiIl , OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 , OoiloolOiOIoIOolLiOl0OlOiOli0oOOl , OillLliLoolOIiiiILoOILOIloo000iLI , OlLOLoI0iIOLloliOllILlOoIiioOli0L , Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l , O0Loo0iiI0OlLOlOIiILOooOOlIoioOli , OoOi0O0oOoL0looLo0IoOllOOILiLooLl , OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO , OLlOiiLlLoolliOiO0i0lOloio0L0oL00 , OilOI0i0lloo0Lll000I0OIoIOI0lioiO , OlooiiLooL0L00oIIiioLloiIolOoOlLo , OLo0LOlILllLILOIiiiL0LIlLIoLlO0II , OiiOioOIO00LOOLilooiooo0olO0illo0 , OLl0LoLoii00oiOOoilollii000iIOlOI , OLlil0000Oiil0IOOLiloIlliOoLLol0L , OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI , OO0OOILiO000LOILL0OllLi0l0oliLOo0 , OLiLllIIIlo0llILiLloLOoooOLOilI0l , Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl , OiL0IiiliiioOOLliLiiLILlIOloOLL0L , OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi , OllLOLiIilI0oili000OiLilLioIOoIl0 , OOooI0loOL0iiOIoOili0OOOLLiiIiLOl , OLIIiIIIOILl0loi0lO0IiOoolLIloi00 , OoOillIILLoLoOioLloli0OLILlIOOoLo , OlOlO00LLloOiOolOiOLOIiloLil0L0LI , OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO , OlOLIILoL0ll0oooOo0OIoLoOoiLIolol , OIlLOILiLLo0ol0OLlI0IILilILLLlILO , O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i , Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL , OOiIlillllLOI0oOOoILlol0ILoIoOLil , OOIiO0olO0OLlo0liIoiOioiIO00oOIiL , O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 , OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l , OlolLlliLo0O0l0lOOolL0ioI0O0Li00l , Oo0oI0oLOLlloloiiLIIol0LilOlOIliI , OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo , OoiLlL0oiiIloLOoloIL0oLii00IIIoII , Oo0LLillol0loLIo0iOl0oOLlIOlILoIO , OOllOo00o0IlooI0l0io0O00l0OIoiILO , OOiiILlloiOoI0OlilIOoiiLOOLol0IoI , OiiLOILl0iLi0L0ilIIoooLLIoliIIIlO , OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI , OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII , OOLOoolOi0LIo0olO0loLllIlllIiiIiI , OOOLiLOilooIi0Iio00ilILoLIILOoOoI , OL0O0IIio0loL0L0Il0li0i00lliIoOOI , OLLOooI0ILL00ILloiliILLLiioooLliI , OILoli0OIOIIOI0OiliOo0i0OLoliOOiI , O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI , OilOOioILlOIIOL0iioIOIi0oloooOoLl, OOL0o0i0Llo0IiiLlO00oliOILLI00Ool , OI00OiLolooiIIiiILoIliO0O0loolIlI , OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo , OIIOLLOIlOlLoi0oiOioLilOiioiiliLO , OIloLiiOL00oilLo0iiILoOOll0lIlIlO , Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII , O0oill0llILOilo0i0LIoOLIoolL0Il0o , OlliILlLOilOl0LO0O0OilooiIIiOi0Ll , OOLoL0looIOoioIoOooIoLIiIiLiLoiOl , OIoIooIolOilIOlooOlOIIOoilLioOIIO , OiL0LolLLIOlliloII00llOil0oIlOiIo , O0llIOIliLOO0iiOoO0OO0lIOloLoII0I , OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL , OilOIloOO0LiLoIL0IIILoIi0Loilll0I , Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 , OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O , OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO , OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 , OlOI0loIIIlOi0OOloOioOIo0L00iOiOi , OO0LlIOOoILoolO0LlO0O0liOIl0OiOil , OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL , OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 , OiooiLLioLLL0lII00ol0oIOllLlOiLlL , OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi , O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 , Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO , O0i0IiOL0liOOoLoOiioLOiIIioolOlLI , OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o , OilLIO0lI0LO0LolOOilILl0oiIlolOlo , OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O , OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL , OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 , OlIIIILlOLoIIio0lIloiiLOIOoliL0IO , OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO , OIoliiOo0i000ooilOOLOiil0LlLiOoLo , Oo00OlooOo0io0OoIloiioLiOlL0llio0 , OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL , OOoOoILioOoIlIoLliOLOOi0io0IlLolo , OiLllooo0Li0lioiolLi0ILIoLOliil0I , OlioIL00LLooOiOiOi0liiLI0OOLLI0lO , OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl , OlIlI0o0I0ILOloiOioI0i0IiIliLil00 , OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo , OLL0OiLILloil0IoOlLIIloLIiIlllLil , OILI0LLillilOlllLil0ioLoIiliOoLLo , OiIOlO00OOiiOlOloOOIl0IIoL00IOliL , OoIloII0oLiOLOLIllOL0iOoooOliOIii , Ol0iOoOil0il0LilI0Io0IIooll0i0I0o , OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL , OO0liOO0iOOIioool0OoLliiiI0l0ilOo , OiIOLi00lOILlOOL0oLLloL0io0LoIoOL , OLo0oiiL0ooIliO0I0illLoILiiIoIoOI , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , OOooLlloIiioOOO0LLILl0liiillLILol , OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI , OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 , OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol , OloliIooiiLI0IIlOiL0LLlioILLllL0L , O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO , OioILlIiO0000OoolooO00loIOIloLIoI , OLOl0000OLooLIIo0lIOIOI0lILioolOl , OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII , OoIolLlOIIoIoi00lloLlIoI0lo0iILol , OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI , OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo , OOIIloOlOILliIOILOIOiIlooIOOIL0oO , OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io , OiLOo0loOI00OL0Ooio0OIIlOLiooLOII , OlLilll0ilOLI0IIoO0li0l0OlO00oLIO , O0liLooiLliIoLOllliIlo0ILo0I0oOOl , O0i00oOl00OoIIOIil0LLOi0looIOIL00 , OOLIiil0IlIllLollIl0LIilliOI0iolo );
 parameter OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL = 5'd0 ;
 parameter OiIoi0liOllioIL0IilOLIOIOIiILiioI = 5'd2 ;
 parameter OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO = 5'd4 ;
 parameter OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo = 5'd5 ;
 parameter OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo = 5'd6 ;
 parameter OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 = 5'd7 ;
 parameter OllIlooiolLL00OiIIiOO0iOOiIlLLOoi = 5'd8 ;
 parameter OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L = 5'd9 ;
 parameter OoIlLOiLLl0Il0Ili0Lo0ooLloO00oILL = 5'd10 ;
 parameter O0IloLIOl0I0oli0IOIoOO0lOolioolIl = 5'd11 ;
 parameter O0OiiIi0olIo0IIL0O0OIIolIiIOLllO0 = 5'd12 ;
 parameter OILlioiLloo0oIiI0o0ILOIIiO0IoiOil = 5'd14 ;
 parameter O0Il0i0oII0Lil0IooLoIIliOoOI0oiO0 = 5'd16 ;
 parameter O0OlILLoioIIlIilolliIoIiliIoLlLoL = 5'd18 ;
 parameter OlOLi0Il0l0LOOlOIOiooiilIIOO0I0oL = 5'd20 ;
 parameter OiilO0lI0iIIOio0IIiiOoIoioLL00oOO = 5'd22 ;
 input [31:0] OoIolioOL0iLLOLloI00iIILLiiL0Ooil ;
 input [31:0] Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 ;
 output [3:0] OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI ;
 output OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 ;
 output [ 5:0] OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI ;
 output OilOOo00lLiOOoiO0ii0oo0oOliOollii ;
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input [15:0] Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 input [15:0] OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ;
 input [15:0] OoiloolOiOIoIOolLiOl0OlOiOli0oOOl ;
 input [15:0] OillLliLoolOIiiiILoOILOIloo000iLI ;
 input [15:0] OlLOLoI0iIOLloliOllILlOoIiioOli0L ;
 output O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ;
 output [31:0] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 input [31:0] OoOi0O0oOoL0looLo0IoOllOOILiLooLl ;
 input [31:0] OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO ;
 input [31:0] OLlOiiLlLoolliOiO0i0lOloio0L0oL00 ;
 input [31:0] OilOI0i0lloo0Lll000I0OIoIOI0lioiO ;
 input [31:0] OlooiiLooL0L00oIIiioLloiIolOoOlLo ;
 input [31:0] OLo0LOlILllLILOIiiiL0LIlLIoLlO0II ;
 input [31:0] OiiOioOIO00LOOLilooiooo0olO0illo0 ;
 input [31:0] OLl0LoLoii00oiOOoilollii000iIOlOI ;
 input [31:0] OLlil0000Oiil0IOOLiloIlliOoLLol0L ;
 input [31:0] OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI ;
 input [31:0] OO0OOILiO000LOILL0OllLi0l0oliLOo0 ;
 input [31:0] OLiLllIIIlo0llILiLloLOoooOLOilI0l ;
 input [31:0] Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl ;
 input [31:0] OiL0IiiliiioOOLliLiiLILlIOloOLL0L ;
 input [31:0] OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi ;
 input [31:0] OllLOLiIilI0oili000OiLilLioIOoIl0 ;
 input [31:0] OOooI0loOL0iiOIoOili0OOOLLiiIiLOl ;
 input [31:0] OLIIiIIIOILl0loi0lO0IiOoolLIloi00 ;
 input [31:0] OoOillIILLoLoOioLloli0OLILlIOOoLo ;
 input [31:0] OlOlO00LLloOiOolOiOLOIiloLil0L0LI ;
 input [31:0] OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO ;
 input [31:0] OlOLIILoL0ll0oooOo0OIoLoOoiLIolol ;
 input [31:0] OIlLOILiLLo0ol0OLlI0IILilILLLlILO ;
 input [31:0] O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i ;
 input [31:0] Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL ;
 input [31:0] OOiIlillllLOI0oOOoILlol0ILoIoOLil ;
 input [31:0] OOIiO0olO0OLlo0liIoiOioiIO00oOIiL ;
 input [31:0] O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 ;
 input [31:0] OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l ;
 input [31:0] OlolLlliLo0O0l0lOOolL0ioI0O0Li00l ;
 input [31:0] Oo0oI0oLOLlloloiiLIIol0LilOlOIliI ;
 input [31:0] OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo ;
 input [31:0] OoiLlL0oiiIloLOoloIL0oLii00IIIoII ;
 input [31:0] Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ;
 input [31:0] OOllOo00o0IlooI0l0io0O00l0OIoiILO ;
 input [31:0] OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ;
 input OiiLOILl0iLi0L0ilIIoooLLIoliIIIlO ;
 input OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ;
 input [ 3:0] OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 input OOLOoolOi0LIo0olO0loLllIlllIiiIiI ;
 input OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 input [63:0] OLLOooI0ILL00ILloiliILLLiioooLliI ;
 input [ 2:0] OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 input [15:0] O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ;
 output OL0O0IIio0loL0L0Il0li0i00lliIoOOI ;
 input [15:0] OilOOioILlOIIOL0iioIOIi0oloooOoLl;
 input [31:0] OOL0o0i0Llo0IiiLlO00oliOILLI00Ool ;
 input OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 input OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ;
 output [31:0] OIloLiiOL00oilLo0iiILoOOll0lIlIlO ;
 output Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ;
 output O0oill0llILOilo0i0LIoOLIoolL0Il0o ;
 output OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ;
 output OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ;
 output OIoIooIolOilIOlooOlOIIOoilLioOIIO ;
 output OiL0LolLLIOlliloII00llOil0oIlOiIo ;
 output O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ;
 output OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL ;
 input [15:0] OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ;
 input OOooLlloIiioOOO0LLILl0liiillLILol ;
 output [31:0] OilOIloOO0LiLoIL0IIILoIi0Loilll0I ;
 output [31:0] Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ;
 output [31:0] OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ;
 output [63:0] OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ;
 output [ 2:0] OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ;
 output [ 2:0] OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ;
 output [ 2:0] OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ;
 output [ 2:0] OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ;
 output [ 2:0] OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ;
 output [ 2:0] OiooiLLioLLL0lII00ol0oIOllLlOiLlL ;
 output [ 2:0] OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ;
 output [ 2:0] O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ;
 output [ 2:0] Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ;
 output [ 2:0] O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ;
 output [ 2:0] OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ;
 output [ 2:0] OilLIO0lI0LO0LolOOilILl0oiIlolOlo ;
 output [ 2:0] OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ;
 output [ 2:0] OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ;
 output [ 2:0] OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ;
 output [ 2:0] OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ;
 output [ 2:0] OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ;
 output [ 2:0] OIoliiOo0i000ooilOOLOiil0LlLiOoLo ;
 output [ 2:0] Oo00OlooOo0io0OoIloiioLiOlL0llio0 ;
 output [ 2:0] OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ;
 output [ 2:0] OOoOoILioOoIlIoLliOLOOi0io0IlLolo ;
 output [ 2:0] OiLllooo0Li0lioiolLi0ILIoLOliil0I ;
 output [ 2:0] OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ;
 output [ 2:0] OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ;
 output [ 2:0] OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ;
 output [ 2:0] OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ;
 output [ 2:0] OLL0OiLILloil0IoOlLIIloLIiIlllLil ;
 output [ 2:0] OILI0LLillilOlllLil0ioLoIiliOoLLo ;
 output [ 2:0] OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ;
 output [ 2:0] OoIloII0oLiOLOLIllOL0iOoooOliOIii ;
 output [ 2:0] Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ;
 output [ 2:0] OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ;
 output [31:0] OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 output OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 output [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 output [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 output [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 output [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 output [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 output [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 output [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 output [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 output [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 output [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 output [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 output [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 output [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 output [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 output [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 output [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 output O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 output [ 15: 0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 output [ 5: 0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 output [ 15: 0] O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ;
 output [ 15:0] OILIloOoilLIL00IIOoOilLOO0L0iiIOO ;
 output [ 31:0] O0oLLi0Ill00l0lioiLioiooIllloIiIl ;
 output OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 output OOLIiil0IlIllLollIl0LIilliOI0iolo;
 input [3:0] Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L ;
 input [3:0] OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl ;
 reg OliOOOIooO0oILLiLiiilLIlilo0ooL0O ;
 wire O0il0IO0olIoLiOIL0000lo0OoliIL0Ll ;
 wire OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 = O0il0IO0olIoLiOIL0000lo0OoliIL0Ll ;
 reg [31:0] OIloLiiOL00oilLo0iiILoOOll0lIlIlO ;
 wire OL0O0IIio0loL0L0Il0li0i00lliIoOOI ;
 reg [ 5:0] Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ;
 reg O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ;
 wire [ 5:0] OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI = Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ;
 wire OilOOo00lLiOOoiO0ii0oo0oOliOollii = O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ;
 wire [31:0] OilOIloOO0LiLoIL0IIILoIi0Loilll0I ;
 wire [31:0] Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ;
 wire [31:0] OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ;
 wire [63:0] OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ;
 wire [ 2:0] OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ;
 wire [ 2:0] OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ;
 wire [ 2:0] OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ;
 wire [ 2:0] OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ;
 wire [ 2:0] OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ;
 wire [ 2:0] OiooiLLioLLL0lII00ol0oIOllLlOiLlL ;
 wire [ 2:0] OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ;
 wire [ 2:0] O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ;
 wire [ 2:0] Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ;
 wire [ 2:0] O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ;
 wire [ 2:0] OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ;
 wire [ 2:0] OilLIO0lI0LO0LolOOilILl0oiIlolOlo ;
 wire [ 2:0] OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ;
 wire [ 2:0] OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ;
 wire [ 2:0] OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ;
 wire [ 2:0] OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ;
 wire [ 2:0] OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ;
 wire [ 2:0] OIoliiOo0i000ooilOOLOiil0LlLiOoLo ;
 wire [ 2:0] Oo00OlooOo0io0OoIloiioLiOlL0llio0 ;
 wire [ 2:0] OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ;
 wire [ 2:0] OOoOoILioOoIlIoLliOLOOi0io0IlLolo ;
 wire [ 2:0] OiLllooo0Li0lioiolLi0ILIoLOliil0I ;
 wire [ 2:0] OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ;
 wire [ 2:0] OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ;
 wire [ 2:0] OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ;
 wire [ 2:0] OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ;
 wire [ 2:0] OLL0OiLILloil0IoOlLIIloLIiIlllLil ;
 wire [ 2:0] OILI0LLillilOlllLil0ioLoIiliOoLLo ;
 wire [ 2:0] OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ;
 wire [ 2:0] OoIloII0oLiOLOLIllOL0iOoooOliOIii ;
 wire [ 2:0] Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ;
 wire [ 2:0] OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ;
 wire [191:0] O0lOIlooLi0lilOllLlilIo00iOLiOLLo ;
 wire [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 wire [ 5:0] OI0iIoio000lOoOiiiI0Loo0l0I0liioO = O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 reg [31:0] OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 reg [31:0] OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0 ;
 reg OOOll0oL0OOLoi0lIioOo0liiLILLoiiL ;
 reg OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 reg [31:0] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 reg OllII0i0lILiOLIL0OiIIoLoiIl0IoLoI ;
 reg OoILOLi0I0lO0LOI0Illoo0Lo0ilOLLoL ;
 reg OOOLIoiLiLOOLooIoOoioiooIIoliLOlo ;
 reg O0llLOll00OIl0OoLOiOiioIo0O0IolOo ;
 reg OlIiOlLoi0loOiLoLoioiIOIioliiLill ;
 reg OOlL0lLllIOooOI0Ol0L0olliOLO0IlII ;
 reg O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ;
 reg [31:0] OoloOOilIOLlIlIII0oIL0IOllO0oLi0o ;
 reg [31:0] O0OoOIloiOI0oOil0LlIl0oil0iLOOiLL ;
 reg [31:0] OlLO0OLOOiLioiL0ILLllii0OlIiOOIo0 ;
 reg [31:0] O0OIlIIlo00lILOO0iOiIILOOI0OI0oOi ;
 reg [31:0] O0i0lIILioOLiLOIiIO00loi0iLOloLLL ;
 reg [31:0] OoLl0IIIo0IollLoILOLlOIiioIIi0iIo ;
 reg [31:0] OIoIi0IlLoooi0iILio0lILiIOL0oLOol ;
 reg [31:0] OIlooiLoolLOlLiOLioooILlolIlIlIoi ;
 reg [31:0] OiloOOiiooL0o0OIOOiiL0Iii0Lii0LLi ;
 reg [31:0] O0O0Il000ILILl0iIOIOOIi00OilLLLoi ;
 reg [31:0] OLoi0olioL0OLoILii0iO00IlOOLI00l0 ;
 reg [31:0] OOlILI0loI0illoollOiIIOl0iii0oIIi ;
 reg [31:0] OiL0iLlILIoiO0lLioo0ololOiILIIoOl ;
 reg [31:0] OlllolOIO000iLIo0I0LoLoOLL0IlLl0O ;
 reg [31:0] OIIOLlIiiOoLOLLoLOOO0OOoOoOLIOool ;
 reg [31:0] OOoLoiLILiiOi0OoO0olOoOoioo0lLoLl ;
 reg [31:0] OLiLOi0l0li0loOLOIolIOIIOiLlilolI ;
 reg [31:0] OlLIiII0LOiOOo0OoloIILoOIoIOi0O00 ;
 reg [31:0] O0OLOILIl0iOLLOoL0LIOIooloLOLo0ii ;
 reg [31:0] OLLOi0ioLIIiliILllOIIioOl0OLilili ;
 reg [31:0] OLi0IOOoOL00iloIi0i0lLioLiIoioOoo ;
 reg [31:0] OIoO0O0OIiIIi00OLLl0olOIOiiIIl0IO ;
 reg [31:0] OoIlOlOiL0ollilOlli00LlIOlioLi0l0 ;
 reg [31:0] OOllii0LlOLLLoLOIOOiiIO0LlIoooOIL ;
 reg [31:0] OoilOILoi0lOli00o0lol0ILilOolil0l ;
 reg [31:0] OLOLOILIoOlIiL0iLOooilloILI0OiLlo ;
 reg [31:0] O0ooio00O00Ii0l0iill0iLLOLLOOOIIo ;
 reg [31:0] OoOOo0iiI0iLoIooI0OIOOiLO0IooOILO ;
 reg [31:0] OoIOL0IiLi0i0Loi0llllioOoiIoOLLIo ;
 reg [31:0] OliLLl0OlLIiOlIIiLlLlooO0LoiLiooO ;
 reg [31:0] OioioLOliOLI0IOlLOolII0L0oi0oIiLO ;
 reg [31:0] O0l0LioII0IlliOlIIi0IlI00IoOOoiOo ;
 wire [15:0] OILIloOoilLIL00IIOoOilLOO0L0iiIOO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:112+64];
 wire [15:0] O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 96+64];
 wire [31:0] O0oLLi0Ill00l0lioiLioiooIllloIiIl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 64+64];
 wire [15:0] Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:112+64];
 wire [31:0] OlO0Oo0looiIoIiL0liIllLLLL0o00i0L = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 80+64];
 wire [31:0] O0o0loiLIOlLoi0iOIolL0LoOILoilLLl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:96+64] ;
 wire [15:0] Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64:80+64] ;
 wire [15:0] OiO0oiLLillil0LLLOLo0OoiiOLLIILiI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 79+64:64+64] ;
 wire [15:0] OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:112+64];
 wire [15:0] OOioILiL0oiO0OIlLLOLLi0O0oOOIlIlI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 96+64];
 wire [15:0] OOiLiOlo0ioloILilO0IlILL0o0iiLiOI = 16'd81 ;
 reg [31:0] Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 reg [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 reg OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 reg [15:0] OLlOlo0lOII0I0i0l0lOiOl0L0iioO0Io ;
 reg [15:0] O0IIOiLIOiIi0Ol0000ilIill0II0OilI ;
 wire [11:0] OlI0LilLLoO0OiiLioLoIIILooLIlILOi ;
 wire [ 3:0] Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ;
 reg [11:0] OOOi0LIiLLOLIoliiOlolloOli0oLLioi ;
 assign OlI0LilLLoO0OiiLioLoIIILooLIlILOi = O0IIOiLIOiIi0Ol0000ilIill0II0OilI[15:4] ;
 assign Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 = O0IIOiLIOiIi0Ol0000ilIill0II0OilI[ 3:0] ;
 wire [3:0] OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI = O0IIOiLIOiIi0Ol0000ilIill0II0OilI[ 3:0] ;
 reg [15:0] OILLIiOoiIOiIil0OLOLLiIIllIlOLilI ;
 reg [15:0] OLIiiio00OOiooIiolIO0ooLl0OlIoloI ;
 reg [15:0] OliiLIIliIO0OIloloLiiI0ilOILLILOI ;
 reg [15:0] OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo ;
 reg [15:0] OLOlIOIOOlLOII0OLL0oiL0I0O0IilloL ;
 wire [11:0] O0oioIoloolL0oiioLILllioiO0oliIOl ;
 wire [ 3:0] Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 assign O0oioIoloolL0oiioLILllioiO0oliIOl = OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo[15:4] ;
 assign Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi = OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo[ 3:0] ;
 reg [11:0] OLIo0LL0IiLIOliLL00I0LO00IllOOllo ;
 reg [15:0] Oi0ILolLOL0li0iLIolliilIlLlloolO0 ;
 wire OIlii0Io00iIi0iIOilOOoollO0iI0lol = OOOLiLOilooIi0Iio00ilILoLIILOoOoI && OL0O0IIio0loL0L0Il0li0i00lliIoOOI ;
 reg OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ;
 assign OL0O0IIio0loL0L0Il0li0i00lliIoOOI = 1'b1 ;
 reg Oiiii0oOiIIl0i00oIOoioo0OiolIooLO ;
 reg OolLol00lliiIOoololoo00lIlIoo0O0I ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oiiii0oOiIIl0i00oIOoioo0OiolIooLO <= 1'd0 ;
 OolLol00lliiIOoololoo00lIlIoo0O0I <= 1'd0 ;
 end
 else begin
 Oiiii0oOiIIl0i00oIOoioo0OiolIooLO <= (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00==OoiloolOiOIoIOolLiOl0OlOiOli0oOOl)|| (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00==OlLOLoI0iIOLloliOllILlOoIiioOli0L);
 OolLol00lliiIOoololoo00lIlIoo0O0I <= (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00==OillLliLoolOIiiiILoOILOIloo000iLI);
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI <= 5'd0 ;
 end
 else begin
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI <= (&OOllOo00o0IlooI0l0io0O00l0OIoiILO) ;
 end
 end
 reg [ 4:0] OOLIiil0IlIllLollIl0LIilliOI0iolo ;
 reg [ 4:0] OL0II0lIOioLIIOLlLILoioOiOLLlLLLL ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLIiil0IlIllLollIl0LIilliOI0iolo <= 5'd0 ;
 end
 else if ( (OiiLOILl0iLi0L0ilIIoooLLIoliIIIlO&&~Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII)||OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) begin
 OOLIiil0IlIllLollIl0LIilliOI0iolo <= 5'd0 ;
 end
 else begin
 OOLIiil0IlIllLollIl0LIilliOI0iolo <= OL0II0lIOioLIIOLlLILoioOiOLLlLLLL ;
 end
 end
 wire Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL );
 wire OlliILlLOilOl0LO0O0OilooiIIiOi0Ll = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OiIoi0liOllioIL0IilOLIOIOIiILiioI );
 wire O0LO0iloLil0LI0IOiOolIoioLOOIOLiO = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO );
 wire OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo );
 wire OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo );
 wire OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 );
 wire OOIIIOLL0O000ioLliOIoOii0LiI0lOoo = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OllIlooiolLL00OiIIiOO0iOOiIlLLOoi );
 wire OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L );
 wire Oo0LiLOLOIi0lLoOlLLiIoo00lLlloOlO = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OoIlLOiLLl0Il0Ili0Lo0ooLloO00oILL );
 wire OLIoo0OL0oo0iloLooi0iIIoLLOlIILIL = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== O0IloLIOl0I0oli0IOIoOO0lOolioolIl );
 wire OOLoL0looIOoioIoOooIoLIiIiLiLoiOl = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== O0OiiIi0olIo0IIL0O0OIIolIiIOLllO0 );
 wire OIoIooIolOilIOlooOlOIIOoilLioOIIO = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OILlioiLloo0oIiI0o0ILOIIiO0IoiOil );
 wire O0oill0llILOilo0i0LIoOLIoolL0Il0o = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== O0Il0i0oII0Lil0IooLoIIliOoOI0oiO0 );
 wire OiL0LolLLIOlliloII00llOil0oIlOiIo = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== O0OlILLoioIIlIilolliIoIiliIoLlLoL );
 wire O0llIOIliLOO0iiOoO0OO0lIOloLoII0I = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OlOLi0Il0l0LOOlOIOiooiilIIOO0I0oL );
 wire O0IIOOO0LOOiLiiOill00LllllIOIILo0 = ( OOLIiil0IlIllLollIl0LIilliOI0iolo== OiilO0lI0iIIOio0IIiiOoIoioLL00oOO ) ;
 always@ ( * ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OOLIiil0IlIllLollIl0LIilliOI0iolo;
 case(OOLIiil0IlIllLollIl0LIilliOI0iolo) OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL : begin
 if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI&&OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OI00OiLolooiIIiiILoIliO0O0loolIlI) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = ( Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l>16'd8 ) ? O0OlILLoioIIlIilolliIoIiliIoLlLoL : OlOLi0Il0l0LOOlOIOiooiilIIOO0I0oL ;
 end
 end
 O0OlILLoioIIlIilolliIoIiliIoLlLoL : begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l<=16'd16) ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OlOLi0Il0l0LOOlOIOiooiilIIOO0I0oL ;
 end
 end
 OlOLi0Il0l0LOOlOIOiooiilIIOO0I0oL : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = ( OolIOLOooiLLIllI0LOLIolllLoilolIl>(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8) ) ? OiIoi0liOllioIL0IilOLIOIOIiILiioI : OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L ;
 end
 end
 OiIoi0liOllioIL0IilOLIOIOIiILiioI : begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) begin
 if ( (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && (OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 if ( OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0&&~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ? (OolIOLOooiLLIllI0LOLIolllLoilolIl<= (16'd8+16'd8) ) ? OILlioiLloo0oIiI0o0ILOIIiO0IoiOil : O0OiiIi0olIo0IIL0O0OIIolIiIOLllO0 : OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 else if ((OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiilO0lI0iIIOio0IIiiOoIoioLL00oOO ;
 end
 end
 end
 OLLoIlioLLlLOi0OL0ii0ILlLi0looIlO : begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd6 ) begin
 if ( ( ((Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OillLliLoolOIiiiILoOILOIloo000iLI)&&OolLol00lliiIOoololoo00lIlIoo0O0I) || ( Oiiii0oOiIIl0i00oIOoioo0OiolIooLO&&((Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OoiloolOiOIoIOolLiOl0OlOiOli0oOOl)||(Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OlLOLoI0iIOLloliOllILlOoIiioOli0L)) ) ) && (OlO0Oo0looiIoIiL0liIllLLLL0o00i0L==32'h0000_5902) ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiilO0lI0iIIOio0IIiiOoIoioLL00oOO ;
 end
 end
 end
 OIOLllOoIoi0Loo0l0iLlL0LiiI0LolLo : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) begin
 if ( (Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI<=16'h0001) || ~OliOOOIooO0oILLiLiiilLIlilo0ooL0O ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoIlLOiLLl0Il0Ili0Lo0ooLloO00oILL ;
 end
 else if ( O0o0loiLIOlLoi0iOIolL0LoOILoilLLl<=OO0liOO0iOOIioool0OoLliiiI0l0ilOo ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoIlLOiLLl0Il0Ili0Lo0ooLloO00oILL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo ;
 end
 end
 end
 OoIlLOiLLl0Il0Ili0Lo0ooLloO00oILL : begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi>=(OlI0LilLLoO0OiiLioLoIIILooLIlILOi-1'b1)) ) begin
 if ( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0==4'd0 ) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl==6'd16 ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else if (OolIOLOooiLLIllI0LOLIolllLoilolIl<=(16'd16+16'd8)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = ( (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli&&OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0) ) ? OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L : OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else if ( OolIOLOooiLLIllI0LOLIolllLoilolIl<(16'd16+ OOiLiOlo0ioloILilO0IlILL0o0iiLiOI ) ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = ( (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli&&OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0) ) ? OiIoi0liOllioIL0IilOLIOIOIiILiioI : OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiIoi0liOllioIL0IilOLIOIOIiILiioI ;
 end
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = O0IloLIOl0I0oli0IOIoOO0lOolioolIl ;
 end
 end
 end
 O0IloLIOl0I0oli0IOIoOO0lOolioolIl: begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl==Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else if (OolIOLOooiLLIllI0LOLIolllLoilolIl<=(Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0+16'd8)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = ( (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli&&OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0) ) ? OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L : OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else if ( OolIOLOooiLLIllI0LOLIolllLoilolIl<( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 + OOiLiOlo0ioloILilO0IlILL0o0iiLiOI )) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = ( (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli&&OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0) ) ? OiIoi0liOllioIL0IilOLIOIOIiILiioI : OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiIoi0liOllioIL0IilOLIOIOIiILiioI ;
 end
 end
 end
 OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4 )begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 ;
 end
 end
 OIiOIiiiI0o0OIi0Ll0OOilLoIOIiooI0 : begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) )begin
 if (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl>( 16'd16 + 16'd8 ) ) OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiIoi0liOllioIL0IilOLIOIOIiILiioI ;
 else OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo ;
 end
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OllIlooiolLL00OiIIiOO0iOOiIlLLOoi ;
 end
 end
 end
 OllIlooiolLL00OiIIiOO0iOOiIlLLOoi : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl>( Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi + 16'd8 ) ) OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OiIoi0liOllioIL0IilOLIOIOIiILiioI ;
 else OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OoloOIo0O0OoIOooLi0iIoL0LOolIOoOo ;
 end
 end
 end
 OL00OlIOo0IiIlILlLilOIoilO0Oo0L0L : begin
 if ( (OolIOLOooiLLIllI0LOLIolllLoilolIl==16'd0) || (OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI&&OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0) ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 else begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ? O0Il0i0oII0Lil0IooLoIIliOoOI0oiO0 : OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 O0Il0i0oII0Lil0IooLoIIliOoOI0oiO0 : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 O0OiiIi0olIo0IIL0O0OIIolIiIOLllO0 : begin
 if ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)&&(OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd16)) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OILlioiLloo0oIiI0o0ILOIIiO0IoiOil ;
 end
 end
 OILlioiLloo0oIiI0o0ILOIIiO0IoiOil : begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 end
 OiilO0lI0iIIOio0IIiiOoIoioLL00oOO : begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 default : begin
 OL0II0lIOioLIIOLlLILoioOiOLLlLLLL = OilIOO0oOLIOiLIiOL0lioIIilLoIiIiL ;
 end
 endcase end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 <= 1'd0 ;
 OliOOOIooO0oILLiLiiilLIlilo0ooL0O <= 1'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 <= OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 OliOOOIooO0oILLiLiiilLIlilo0ooL0O <= OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 end
 else if ( O0LO0iloLil0LI0IOiOolIoioLOOIOLiO ) begin
 OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 <= ( ((Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OillLliLoolOIiiiILoOILOIloo000iLI)&&OolLol00lliiIOoololoo00lIlIoo0O0I) || ( Oiiii0oOiIIl0i00oIOoioo0OiolIooLO&&((Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OoiloolOiOIoIOolLiOl0OlOiOli0oOOl)||(Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OlLOLoI0iIOLloliOllILlOoIiioOli0L)) ) ) ;
 OliOOOIooO0oILLiLiiilLIlilo0ooL0O <= (Oll0IOoii0OiilO00OIoL0iLiIiiiOLLO==OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00) ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLlOlo0lOII0I0i0l0lOiOl0L0iioO0Io <= 16'd0 ;
 end
 else if ( ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OLlOlo0lOII0I0i0l0lOiOl0L0iioO0Io <= O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0IIOiLIOiIi0Ol0000ilIill0II0OilI <= 16'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI) begin
 O0IIOiLIOiIi0Ol0000ilIill0II0OilI <= OilOOioILlOIIOL0iioIOIi0oloooOoLl - 16'd22 ;
 end
 else if ( ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 O0IIOiLIOiIi0Ol0000ilIill0II0OilI <= O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo - 16'd22 ;
 end
 end
 reg OlIl0ooIoiLlO0lII0loOOi0IoIILloOO ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlIl0ooIoiLlO0lII0loOOi0IoIILloOO <= 1'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI) begin
 if (OilOOioILlOIIOL0iioIOIi0oloooOoLl==16'd0) begin
 OlIl0ooIoiLlO0lII0loOOi0IoIILloOO <= 1'd1 ;
 /* synthesis translate_off */ $display("%m OilOOioILlOIIOL0iioIOIi0oloooOoLl = %d Error !!!!! \n ", OilOOioILlOIIOL0iioIOIi0oloooOoLl );
 /* synthesis translate_on */ end
 else begin
 OlIl0ooIoiLlO0lII0loOOi0IoIILloOO <= 1'd0 ;
 end
 end
 else begin
 OlIl0ooIoiLlO0lII0loOOi0IoIILloOO <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= 16'd0 ;
 end
 else if ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && ~OI00OiLolooiIIiiILoIliO0O0loolIlI ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= (O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI<=16'd8) ? (OIIOLLOIlOlLoi0oiOioLilOiioiiliLO - OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ) : (OIIOLLOIlOlLoi0oiOioLilOiioiiliLO - O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI - OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII + 16'd8 ) ;
 end
 else if ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OI00OiLolooiIIiiILoIliO0O0loolIlI ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= (OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ) ;
 end
 else if ( Oo0LiLOLOIi0lLoOlLLiIoo00lLlloOlO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd16) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd16 ;
 end
 else if ( OLIoo0OL0oo0iloLooi0iIIoLLOlIILIL && ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if (O0LO0iloLil0LI0IOiOolIoioLOOIOLiO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd6) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd6 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd12) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd12 ;
 end
 else if (OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd4) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd4 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd16 ;
 end
 else if (OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 end
 else if ( OOLoL0looIOoioIoOooIoLIiIiLiLoiOl && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if ( OIoIooIolOilIOlooOlOIIOoilLioOIIO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ( (O0oill0llILOilo0i0LIoOLIoolL0Il0o ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ((OiL0LolLLIOlliloII00llOil0oIlOiIo) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - 16'd8 ;
 end
 else if ((O0llIOIliLOO0iiOoO0OO0lIOloLoII0I) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l) ) begin
 OolIOLOooiLLIllI0LOLIolllLoilolIl <= OolIOLOooiLLIllI0LOLIolllLoilolIl - Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOOi0LIiLLOLIoliiOlolloOli0oLLioi <= 12'd0 ;
 end
 else if ( Oo0LiLOLOIi0lLoOlLLiIoo00lLlloOlO||OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li ) begin
 OOOi0LIiLLOLIoliiOlolloOli0oLLioi <= (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) ? OOOi0LIiLLOLIoliiOlolloOli0oLLioi + 1'd1 : OOOi0LIiLLOLIoliiOlolloOli0oLLioi ;
 end
 else begin
 OOOi0LIiLLOLIoliiOlolloOli0oLLioi <= 12'd0 ;
 end
 end
 reg OIoOolllLOOiliOLL0oOLo0LLloIOOi0l ;
 reg OOoIliOliILLi0IiIlILLo00iLoLiloIl ;
 reg OIIILoOLllIiLloiiIoiiLooiiI00Oii0 ;
 reg OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 ;
 reg OI00liOIoliolOollOLoioOLooloiloI0 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo <= 16'd0 ;
 OLOlIOIOOlLOII0OLL0oiL0I0O0IilloL <= 16'd0 ;
 OIoOolllLOOiliOLL0oOLo0LLloIOOi0l <= 1'd0 ;
 OOoIliOliILLi0IiIlILLo00iLoLiloIl <= 1'd0 ;
 OIIILoOLllIiLloiiIoiiLooiiI00Oii0 <= 1'd0 ;
 end
 else if ( OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4) ) begin
 OiiilOIlOoI0o0iLOIIl0OIOOlioILlLo <= OOioILiL0oiO0OIlLLOLLi0O0oOOIlIlI ;
 OLOlIOIOOlLOII0OLL0oiL0I0O0IilloL <= OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL ;
 OIoOolllLOOiliOLL0oOLo0LLloIOOi0l <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2439) ;
 OOoIliOliILLi0IiIlILLo00iLoLiloIl <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2433) ;
 OIIILoOLllIiLloiiIoiiLooiiI00Oii0 <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2434) ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 <= 1'd0 ;
 OI00liOIoliolOollOLoioOLooloiloI0 <= 1'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 <= 1'd0 ;
 OI00liOIoliolOollOLoioOLooloiloI0 <= 1'd0 ;
 end
 else if ( OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4) ) begin
 OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2433) ? 1'd1 : OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 ;
 OI00liOIoliolOollOLoioOLooloiloI0 <= (OolOoLOOliLoIIO0lo0ilLiiLooLoo0LL==16'h2434) ? 1'd1 : OI00liOIoliolOollOLoioOLooloiloI0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OILLIiOoiIOiIil0OLOLLiIIllIlOLilI <= 16'd0 ;
 OLIiiio00OOiooIiolIO0ooLl0OlIoloI <= 16'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) ) begin
 OILLIiOoiIOiIil0OLOLLiIIllIlOLilI <= Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI ;
 OLIiiio00OOiooIiolIO0ooLl0OlIoloI <= OiO0oiLLillil0LLLOLo0OoiiOLLIILiI ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OliiLIIliIO0OIloloLiiI0ilOILLILOI <= 16'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OliiLIIliIO0OIloloLiiI0ilOILLILOI <= 16'd0 ;
 end
 else if ( OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4 ) ) begin
 OliiLIIliIO0OIloloLiiI0ilOILLILOI <= OliiLIIliIO0OIloloLiiI0ilOILLILOI + 1'd1 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI && OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII<=3'd2) ? 6'd6 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII<=3'd2) ? 1'd1 : 1'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OI00OiLolooiIIiiILoIliO0O0loolIlI && OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l>16'd8) ? ( (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII==3'd0) ? 6'd8 : 6'd0 ) : ((Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[3:0]+OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII)>4'd8) ? 6'd0 : Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[3:0] ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l>16'd8) ? ( (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII==3'd0) ? 1'd1 : 1'd0 ) : ((Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[3:0]+OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII)>4'd8) ? 1'd0 : 1'd1 ;
 end
 else if (OiL0LolLLIOlliloII00llOil0oIlOiIo) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l<=16'd16) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]))) ? Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] - 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= (OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]))) ? 1'd1 : 1'd0;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I && ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8)))&&(OolIOLOooiLLIllI0LOLIolllLoilolIl>(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8))) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((OIlii0Io00iIi0iIOilOOoollO0iI0lol || (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8)))&&(OolIOLOooiLLIllI0LOLIolllLoilolIl>(Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0]+6'd8))) ? 1'd1 : 1'd0 ;
 end
 else if (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I && OIlii0Io00iIi0iIOilOOoollO0iI0lol ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) begin
 if ( OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4 ) ) begin
 if ( (OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0&&O0Loo0iiI0OlLOlOIiILOooOOlIoioOli&&~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ) &&(OolIOLOooiLLIllI0LOLIolllLoilolIl<=(16'd8+16'd8) )) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl[5:0])||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? (OolIOLOooiLLIllI0LOLIolllLoilolIl[5:0]-6'd8) : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl[5:0])||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 end
 else if ((OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd14)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd6 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd14)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (O0LO0iloLil0LI0IOiOolIoioLOOIOLiO) begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd6 ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd18)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd10))) ? 6'd12 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd18)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd10))) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd6 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) begin
 if ( (O0o0loiLIOlLoi0iOIolL0LoOILoilLLl<=OO0liOO0iOOIioool0OoLliiiI0l0ilOo) || (Oo0LlOiOLOl0ooooo0iLOIlo0LILL0iOI<=16'h0001) || ~OliOOOIooO0oILLiLiiilLIlilo0ooL0O ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd28)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20))) ? 6'd16 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd28)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20))) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd4 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd12 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if ( Oo0LiLOLOIi0lLoOlLLiIoo00lLlloOlO ) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi>=(OlI0LilLLoO0OiiLioLoIIILooLIlILOi-1'b1)) ) begin
 if ( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0==4'd0 ) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl<=(16'd16+16'd8)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd24)|| OIlii0Io00iIi0iIOilOOoollO0iI0lol ) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd24)|| OIlii0Io00iIi0iIOilOOoollO0iI0lol ) ? 1'd1 : 1'd0 ;
 end
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd16+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0)))) ? Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd16+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0)))) ? 1'd1 : 1'd0 ;
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? 6'd0 : 6'd16 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? 1'd0 : 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OLIoo0OL0oo0iloLooi0iIIoLLOlIILIL) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ) begin
 if (OolIOLOooiLLIllI0LOLIolllLoilolIl<=( Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 +16'd8)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))|| OIlii0Io00iIi0iIOilOOoollO0iI0lol ) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd8+Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0))|| OIlii0Io00iIi0iIOilOOoollO0iI0lol ) ? 1'd1 : 1'd0 ;
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol && ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8)>= Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oili0OoiliOi0LLoLliiIiIlOiOLOLiL0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OLiLI0Oll0oioO0I0OlI0iOL0LoOlo0iI) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd4 )begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12))) ? 6'd16 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)||(OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12))) ? 1'd1 : 1'd0 ;
 end
 else if ( OIlii0Io00iIi0iIOilOOoollO0iI0lol ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd4 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li) begin
 if ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) )begin
 if (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI<OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd4 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd20)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else if ( OolIOLOooiLLIllI0LOLIolllLoilolIl>( 16'd16 + 16'd8 ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd24)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd24)||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else begin
 if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd16+Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol && ((O0IOooLliOlIllOliILoolIIoIiO0Ilol-6'd8 )>= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol&&(O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? 6'd0 : 6'd16 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? 1'd0 : 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo ) begin
 if ( O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi)begin
 if (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) begin
 if ( OolIOLOooiLLIllI0LOLIolllLoilolIl>( Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi + 16'd8 ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi+16'd8) )||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd8 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi+16'd8) )||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd4+Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi))||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 6'd4 : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(6'd4+Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi))||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 end
 else if ( OIlii0Io00iIi0iIOilOOoollO0iI0lol&& ( (O0IOooLliOlIllOliILoolIIoIiO0Ilol+6'd8) >= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ) ) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else if (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 else if ( OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) begin
 if ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8)&&(OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd16)) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(OolIOLOooiLLIllI0LOLIolllLoilolIl))||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? (OolIOLOooiLLIllI0LOLIolllLoilolIl[5:0]-6'd8) : 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=(OolIOLOooiLLIllI0LOLIolllLoilolIl))||OIlii0Io00iIi0iIOilOOoollO0iI0lol) ? 1'd1 : 1'd0 ;
 end
 else if (OIlii0Io00iIi0iIOilOOoollO0iI0lol) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else if ((O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16)&&O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI) begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd8 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd1 ;
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 else begin
 Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl <= 6'd0 ;
 O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI <= 1'd0 ;
 end
 end
 wire [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 wire [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 reg [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 wire [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 wire [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 reg [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 reg [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 reg [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 reg [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 reg [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 reg [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 reg [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 reg [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 reg [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 reg [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 reg [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 reg O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol <= 32'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) ) begin
 OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol <= {O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[7:0],O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[15:8],O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[23:16],O0o0loiLIOlLoi0iOIolL0LoOILoilLLl[31:24]} ;
 end
 end
 wire [127: 0] OILiOOlOoOl0OiO0OlOoOliIILlliioOl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 64] ;
 wire [ 47: 0] OIIooioLOLO0OIiOiiiooOOIOI0OollII = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:80+64] ;
 wire [ 71: 0] OIlIOllOoilOIlI0OLLoL0l00l0ilooIi = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 79+64: 8+64] ;
 wire [ 7: 0] OiLOLi0io00oIo00Io0lLlLIL0lioiI00 = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 7+64: 64] ;
 wire [ 63: 0] OOILIooliL0iOIOlilO0OiLlLoLIiLOil = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:64+64] ;
 wire [ 31: 0] OOIliIiiiilolLLLLLoi0IlLoilIIOiII = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64:32+64] ;
 wire [ 63: 0] Oo0OioiiiiIiloIIL0ILILoliiO0iooOL = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 64+64] ;
 wire [ 31: 0] OiILllOLOIIl00ooOllolL0OiIIIIOlL0 = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64: 32+64] ;
 wire [ 31: 0] OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 31+64: 64] ;
 wire [ 31: 0] OlooLooOLllollooO0LLIIOilii0o0OlO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 96+64] ;
 wire [ 63: 0] Ol0oii0iIi0Ioo0loOil0000LooOL0OOl = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 32+64] ;
 wire [ 63: 0] OOIOIOIOooiooiilLoOIoL0olL0O0o0Il = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 64+64] ;
 wire [ 31: 0] O0OLLl000lO0LIi0o00iolO0ILoIlOi0O = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64: 32+64] ;
 wire [ 31: 0] OilOOoIIOl0liLOilL0o0LiliIioOLOiI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 31+64: 64] ;
 wire [ 31: 0] OolOIilLOLOLLLiIoOlloool0lolooiO0 = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 96+64] ;
 wire [ 31: 0] OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 64+64] ;
 assign OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI = {8'h53,8'h51,8'h00} ;
 assign OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 = 8'h31 ;
 assign OloliIooiiLI0IIlOiL0LLlioILLllL0L = 8'h30 ;
 assign O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO = 32'd0 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OioILlIiO0000OoolooO00loIOIloLIoI <= 176'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OioILlIiO0000OoolooO00loIOIloLIoI <= 176'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OioILlIiO0000OoolooO00loIOIloLIoI[175:48] <= OILiOOlOoOl0OiO0OlOoOliIILlliioOl ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd1) ) begin
 OioILlIiO0000OoolooO00loIOIloLIoI[47: 0] <= OIIooioLOLO0OIiOiiiooOOIOI0OollII ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl <= 72'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl <= 72'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd1) ) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl[71:64] <= OiLOLi0io00oIo00Io0lLlLIL0lioiI00 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd2) ) begin
 OLOl0000OLooLIIo0lIOIOI0lILioolOl[63: 0] <= OOILIooliL0iOIOlilO0OiLlLoLIiLOil ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIoOolllLOOiliOLL0oOLo0LLloIOOi0l) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd2) ) begin
 OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII[31: 0] <= {OOIliIiiiilolLLLLLoi0IlLoilIIOiII[7:0],OOIliIiiiilolLLLLLoi0IlLoilIIOiII[15:8],OOIliIiiiilolLLLLLoi0IlLoilIIOiII[23:16],OOIliIiiiilolLLLLLoi0IlLoilIIOiII[31:24]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OoIolLlOIIoIoi00lloLlIoI0lo0iILol <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OoIolLlOIIoIoi00lloLlIoI0lo0iILol[63:0]) ) begin
 OoIolLlOIIoIoi00lloLlIoI0lo0iILol <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OoIolLlOIIoIoi00lloLlIoI0lo0iILol[63: 0] <= {Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[7:0],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[15:8],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[23:16],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[31:24],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[39:32],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[47:40],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[55:48],Oo0OioiiiiIiloIIL0ILILoliiO0iooOL[63:56]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI[31: 0] <= { OiILllOLOIIl00ooOllolL0OiIIIIOlL0[7:0],OiILllOLOIIl00ooOllolL0OiIIIIOlL0[15:8],OiILllOLOIIl00ooOllolL0OiIIIIOlL0[23:16],OiILllOLOIIl00ooOllolL0OiIIIIOlL0[31:24] } ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[63:0]) ) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[31: 0] <= { OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[7:0],OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[15:8],OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[23:16],OoO0lOOLiIl0II00oOlOLo0Oo0Loo0Oll[31:24] } ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) ) begin
 OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[63: 32] <= { OlooLooOLllollooO0LLIIOilii0o0OlO[7:0],OlooLooOLllollooO0LLIIOilii0o0OlO[15:8],OlooLooOLllollooO0LLIIOilii0o0OlO[23:16],OlooLooOLllollooO0LLIIOilii0o0OlO[31:24] } ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOIIloOlOILliIOILOIOiIlooIOOIL0oO <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OOIIloOlOILliIOILOIOiIlooIOOIL0oO[63:0]) ) begin
 OOIIloOlOILliIOILOIOiIlooIOOIL0oO <= 'd0 ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OOoIliOliILLi0IiIlILLo00iLoLiloIl) ) begin
 OOIIloOlOILliIOILOIOiIlooIOOIL0oO[63: 0] <= {Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[7:0],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[15:8],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[23:16],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[31:24],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[39:32],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[47:40],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[55:48],Ol0oii0iIi0Ioo0loOil0000LooOL0OOl[63:56]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO || (&OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io[63:0]) ) begin
 OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io[63: 0] <= {OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[7:0],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[15:8],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[23:16],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[31:24],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[39:32],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[47:40],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[55:48],OOIOIOIOooiooiilLoOIoL0olL0O0o0Il[63:56]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiLOo0loOI00OL0Ooio0OIIlOLiooLOII <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 OiLOo0loOI00OL0Ooio0OIIlOLiooLOII <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OiLOo0loOI00OL0Ooio0OIIlOLiooLOII[31: 0] <= {O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[7:0],O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[15:8],O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[23:16],O0OLLl000lO0LIi0o00iolO0ILoIlOi0O[31:24]} ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO <= 64'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO ) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO <= 'd0 ;
 end
 else if ( OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi==12'd0) ) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[31: 0] <= {OilOOoIIOl0liLOilL0o0LiliIioOLOiI[7:0],OilOOoIIOl0liLOilL0o0LiliIioOLOiI[15:8],OilOOoIIOl0liLOilL0o0LiliIioOLOiI[23:16],OilOOoIIOl0liLOilL0o0LiliIioOLOiI[31:24] } ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) ) begin
 OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[63: 0] <= ((&OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[31: 0])&&(&OolOIilLOLOLLLiIoOlloool0lolooiO0[31:0])) ? 64'd0 : { {OolOIilLOLOLLLiIoOlloool0lolooiO0[7:0],OolOIilLOLOLLLiIoOlloool0lolooiO0[15:8],OolOIilLOLOLLLiIoOlloool0lolooiO0[23:16],OolOIilLOLOLLLiIoOlloool0lolooiO0[31:24] } , OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[31:0] } ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0liLooiLliIoLOllliIlo0ILo0I0oOOl <= 32'd0 ;
 end
 else if (OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO) begin
 O0liLooiLliIoLOllliIlo0ILo0I0oOOl <= 'd0 ;
 end
 else if ( OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (OIIILoOLllIiLloiiIoiiLooiiI00Oii0) ) begin
 O0liLooiLliIoLOllliIlo0ILo0I0oOOl[31: 0] <= {OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[7:0],OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[15:8],OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[23:16],OlLLLoIIoLLiO0i00LoIlOIOIii0I0IiO[31:24]} ;
 end
 end
 reg OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= 32'd0 ;
 OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl <= 1'd0 ;
 end
 else begin
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0) 32'h0000_0001: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO) ;
 32'h0000_0002: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLlOiiLlLoolliOiO0i0lOloio0L0oL00) ;
 32'h0000_0004: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OilOI0i0lloo0Lll000I0OIoIOI0lioiO) ;
 32'h0000_0008: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlooiiLooL0L00oIIiioLloiIolOoOlLo) ;
 32'h0000_0010: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLo0LOlILllLILOIiiiL0LIlLIoLlO0II) ;
 32'h0000_0020: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OiiOioOIO00LOOLilooiooo0olO0illo0) ;
 32'h0000_0040: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLl0LoLoii00oiOOoilollii000iIOlOI) ;
 32'h0000_0080: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLlil0000Oiil0IOOLiloIlliOoLLol0L) ;
 32'h0000_0100: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI) ;
 32'h0000_0200: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OO0OOILiO000LOILL0OllLi0l0oliLOo0) ;
 32'h0000_0400: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLiLllIIIlo0llILiLloLOoooOLOilI0l) ;
 32'h0000_0800: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl) ;
 32'h0000_1000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OiL0IiiliiioOOLliLiiLILlIOloOLL0L) ;
 32'h0000_2000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi) ;
 32'h0000_4000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OllLOLiIilI0oili000OiLilLioIOoIl0) ;
 32'h0000_8000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOooI0loOL0iiOIoOili0OOOLLiiIiLOl) ;
 32'h0001_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLIIiIIIOILl0loi0lO0IiOoolLIloi00) ;
 32'h0002_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OoOillIILLoLoOioLloli0OLILlIOOoLo) ;
 32'h0004_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlOlO00LLloOiOolOiOLOIiloLil0L0LI) ;
 32'h0008_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO) ;
 32'h0010_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlOLIILoL0ll0oooOo0OIoLoOoiLIolol) ;
 32'h0020_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OIlLOILiLLo0ol0OLlI0IILilILLLlILO) ;
 32'h0040_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i) ;
 32'h0080_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL) ;
 32'h0100_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOiIlillllLOI0oOOoILlol0ILoIoOLil) ;
 32'h0200_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOIiO0olO0OLlo0liIoiOioiIO00oOIiL) ;
 32'h0400_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0) ;
 32'h0800_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l) ;
 32'h1000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlolLlliLo0O0l0lOOolL0ioI0O0Li00l) ;
 32'h2000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (Oo0oI0oLOLlloloiiLIIol0LilOlOIliI) ;
 32'h4000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo) ;
 32'h8000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OoiLlL0oiiIloLOoloIL0oLii00IIIoII) ;
 default : Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 endcase OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 ;
 end
 end
 reg Oo0iilo0l0ooiililOoLOOL000LLl0OOo ;
 reg [31:0] O0iLolooLLoLIiooi0IlllI0oOll00loO ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0iLolooLLoLIiooi0IlllI0oOll00loO <= 32'd0 ;
 Oo0iilo0l0ooiililOoLOOL000LLl0OOo <= 1'd0 ;
 end
 else begin
 case (OoOi0O0oOoL0looLo0IoOllOOILiLooLl) 32'h0000_0001: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO) ;
 32'h0000_0002: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLlOiiLlLoolliOiO0i0lOloio0L0oL00) ;
 32'h0000_0004: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OilOI0i0lloo0Lll000I0OIoIOI0lioiO) ;
 32'h0000_0008: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OlooiiLooL0L00oIIiioLloiIolOoOlLo) ;
 32'h0000_0010: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLo0LOlILllLILOIiiiL0LIlLIoLlO0II) ;
 32'h0000_0020: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OiiOioOIO00LOOLilooiooo0olO0illo0) ;
 32'h0000_0040: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLl0LoLoii00oiOOoilollii000iIOlOI) ;
 32'h0000_0080: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLlil0000Oiil0IOOLiloIlliOoLLol0L) ;
 32'h0000_0100: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI) ;
 32'h0000_0200: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OO0OOILiO000LOILL0OllLi0l0oliLOo0) ;
 32'h0000_0400: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLiLllIIIlo0llILiLloLOoooOLOilI0l) ;
 32'h0000_0800: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl) ;
 32'h0000_1000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OiL0IiiliiioOOLliLiiLILlIOloOLL0L) ;
 32'h0000_2000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi) ;
 32'h0000_4000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OllLOLiIilI0oili000OiLilLioIOoIl0) ;
 32'h0000_8000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OOooI0loOL0iiOIoOili0OOOLLiiIiLOl) ;
 32'h0001_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OLIIiIIIOILl0loi0lO0IiOoolLIloi00) ;
 32'h0002_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OoOillIILLoLoOioLloli0OLILlIOOoLo) ;
 32'h0004_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OlOlO00LLloOiOolOiOLOIiloLil0L0LI) ;
 32'h0008_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO) ;
 32'h0010_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OlOLIILoL0ll0oooOo0OIoLoOoiLIolol) ;
 32'h0020_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OIlLOILiLLo0ol0OLlI0IILilILLLlILO) ;
 32'h0040_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i) ;
 32'h0080_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL) ;
 32'h0100_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OOiIlillllLOI0oOOoILlol0ILoIoOLil) ;
 32'h0200_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OOIiO0olO0OLlo0liIoiOioiIO00oOIiL) ;
 32'h0400_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0) ;
 32'h0800_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l) ;
 32'h1000_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OlolLlliLo0O0l0lOOolL0ioI0O0Li00l) ;
 32'h2000_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (Oo0oI0oLOLlloloiiLIIol0LilOlOIliI) ;
 32'h4000_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo) ;
 32'h8000_0000: O0iLolooLLoLIiooi0IlllI0oOll00loO <= (OoiLlL0oiiIloLOoloIL0oLii00IIIoII) ;
 default : O0iLolooLLoLIiooi0IlllI0oOll00loO <= O0iLolooLLoLIiooi0IlllI0oOll00loO ;
 endcase Oo0iilo0l0ooiililOoLOOL000LLl0OOo <= |OoOi0O0oOoL0looLo0IoOllOOILiLooLl ;
 end
 end
 reg OiLoLOLiLooLLi0loLlLiooo0LliOiIoL ;
 reg [3:0] OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo <= 32'd0 ;
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= 1'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi || OOOll0oL0OOLoi0lIioOo0liiLILLoiiL ) begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo <= 32'd0 ;
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= 1'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) && OliOOOIooO0oILLiLiiilLIlilo0ooL0O && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ) begin
 if ( O0o0loiLIOlLoi0iOIolL0LoOILoilLLl<=OO0liOO0iOOIioool0OoLliiiI0l0ilOo ) begin
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= 1'd0 ;
 end
 else if (OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo) begin
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= 1'd0 ;
 end
 else if ( (O0o0loiLIOlLoi0iOIolL0LoOILoilLLl<=(OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0+1'd1) ) || (OO0liOO0iOOIioool0OoLliiiI0l0ilOo==32'd0) || (OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl>=OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl) ) begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo <= O0o0loiLIOlLoi0iOIolL0LoOILoilLLl ;
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd1 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= 1'd0 ;
 end
 else begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo <= OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= ((O0o0loiLIOlLoi0iOIolL0LoOILoilLLl-OO0liOO0iOOIioool0OoLliiiI0l0ilOo)>=32'd128 ) ;
 end
 end
 else if (OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl && (OO0liOO0iOOIioool0OoLliiiI0l0ilOo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ) begin
 OO0liOO0iOOIioool0OoLliiiI0l0ilOo <= ((Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO-OO0liOO0iOOIioool0OoLliiiI0l0ilOo)>= 32'd8) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo : Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= ((Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO-OO0liOO0iOOIioool0OoLliiiI0l0ilOo)>=32'd128 ) ;
 end
 else begin
 OiIOLi00lOILlOOL0oLLloL0io0LoIoOL <= 1'd0 ;
 OiLoLOLiLooLLi0loLlLiooo0LliOiIoL <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0 <= 32'd0 ;
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= 4'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi || OOOll0oL0OOLoi0lIioOo0liiLILLoiiL) begin
 OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0 <= 32'd0 ;
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= 4'd0 ;
 end
 else if (Oo0iilo0l0ooiililOoLOOL000LLl0OOo) begin
 if ((O0iLolooLLoLIiooi0IlllI0oOll00loO==(OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0+1'd1)) || (OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl>=OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl) || (OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0==32'd0) ) begin
 OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0 <= (O0iLolooLLoLIiooi0IlllI0oOll00loO) ;
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= 4'd0 ;
 end
 else if (O0iLolooLLoLIiooi0IlllI0oOll00loO>(OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0+1'd1)) begin
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl + 1'd1 ;
 end
 else begin
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= 4'd0 ;
 end
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) && OliOOOIooO0oILLiLiiilLIlilo0ooL0O && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ) begin
 if ( (O0o0loiLIOlLoi0iOIolL0LoOILoilLLl==(OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0+1'd1)) || (OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl>=OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl) || (OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0==32'd0) ) begin
 OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0 <= O0o0loiLIOlLoi0iOIolL0LoOILoilLLl ;
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= 4'd0 ;
 end
 else if (O0o0loiLIOlLoi0iOIolL0LoOILoilLLl>(OIlIiIloLiOOI0OiiLlLL0I00IoioIIo0+1'd1)) begin
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl + 1'd1 ;
 end
 else begin
 OlOLLO0OiOlOLiLOo0lOI0IILLI0iOLIl <= 4'd0 ;
 end
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLo0oiiL0ooIliO0I0illLoILiiIoIoOI <= 32'd0 ;
 OllII0i0lILiOLIL0OiIIoLoiIl0IoLoI <= 1'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OLo0oiiL0ooIliO0I0illLoILiiIoIoOI <= 32'd0 ;
 OllII0i0lILiOLIL0OiIIoLoiIl0IoLoI <= 1'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) && OliOOOIooO0oILLiLiiilLIlilo0ooL0O && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ) begin
 OLo0oiiL0ooIliO0I0illLoILiiIoIoOI <= O0o0loiLIOlLoi0iOIolL0LoOILoilLLl ;
 OllII0i0lILiOLIL0OiIIoLoiIl0IoLoI <= 1'd1 ;
 end
 else begin
 OllII0i0lILiOLIL0OiIIoLoiIl0IoLoI <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OoloOOilIOLlIlIII0oIL0IOllO0oLi0o <= 32'hffff_ffff ;
 O0OoOIloiOI0oOil0LlIl0oil0iLOOiLL <= 32'hffff_ffff ;
 OlLO0OLOOiLioiL0ILLllii0OlIiOOIo0 <= 32'hffff_ffff ;
 O0OIlIIlo00lILOO0iOiIILOOI0OI0oOi <= 32'hffff_ffff ;
 O0i0lIILioOLiLOIiIO00loi0iLOloLLL <= 32'hffff_ffff ;
 OoLl0IIIo0IollLoILOLlOIiioIIi0iIo <= 32'hffff_ffff ;
 OIoIi0IlLoooi0iILio0lILiIOL0oLOol <= 32'hffff_ffff ;
 OIlooiLoolLOlLiOLioooILlolIlIlIoi <= 32'hffff_ffff ;
 OiloOOiiooL0o0OIOOiiL0Iii0Lii0LLi <= 32'hffff_ffff ;
 O0O0Il000ILILl0iIOIOOIi00OilLLLoi <= 32'hffff_ffff ;
 OLoi0olioL0OLoILii0iO00IlOOLI00l0 <= 32'hffff_ffff ;
 OOlILI0loI0illoollOiIIOl0iii0oIIi <= 32'hffff_ffff ;
 OiL0iLlILIoiO0lLioo0ololOiILIIoOl <= 32'hffff_ffff ;
 OlllolOIO000iLIo0I0LoLoOLL0IlLl0O <= 32'hffff_ffff ;
 OIIOLlIiiOoLOLLoLOOO0OOoOoOLIOool <= 32'hffff_ffff ;
 OOoLoiLILiiOi0OoO0olOoOoioo0lLoLl <= 32'hffff_ffff ;
 OLiLOi0l0li0loOLOIolIOIIOiLlilolI <= 32'hffff_ffff ;
 OlLIiII0LOiOOo0OoloIILoOIoIOi0O00 <= 32'hffff_ffff ;
 O0OLOILIl0iOLLOoL0LIOIooloLOLo0ii <= 32'hffff_ffff ;
 OLLOi0ioLIIiliILllOIIioOl0OLilili <= 32'hffff_ffff ;
 OLi0IOOoOL00iloIi0i0lLioLiIoioOoo <= 32'hffff_ffff ;
 OIoO0O0OIiIIi00OLLl0olOIOiiIIl0IO <= 32'hffff_ffff ;
 OoIlOlOiL0ollilOlli00LlIOlioLi0l0 <= 32'hffff_ffff ;
 OOllii0LlOLLLoLOIOOiiIO0LlIoooOIL <= 32'hffff_ffff ;
 OoilOILoi0lOli00o0lol0ILilOolil0l <= 32'hffff_ffff ;
 OLOLOILIoOlIiL0iLOooilloILI0OiLlo <= 32'hffff_ffff ;
 O0ooio00O00Ii0l0iill0iLLOLLOOOIIo <= 32'hffff_ffff ;
 OoOOo0iiI0iLoIooI0OIOOiLO0IooOILO <= 32'hffff_ffff ;
 OoIOL0IiLi0i0Loi0llllioOoiIoOLLIo <= 32'hffff_ffff ;
 OliLLl0OlLIiOlIIiLlLlooO0LoiLiooO <= 32'hffff_ffff ;
 OioioLOliOLI0IOlLOolII0L0oi0oIiLO <= 32'hffff_ffff ;
 O0l0LioII0IlliOlIIi0IlI00IoOOoiOo <= 32'hffff_ffff ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OoloOOilIOLlIlIII0oIL0IOllO0oLi0o <= 32'hffff_ffff ;
 O0OoOIloiOI0oOil0LlIl0oil0iLOOiLL <= 32'hffff_ffff ;
 OlLO0OLOOiLioiL0ILLllii0OlIiOOIo0 <= 32'hffff_ffff ;
 O0OIlIIlo00lILOO0iOiIILOOI0OI0oOi <= 32'hffff_ffff ;
 O0i0lIILioOLiLOIiIO00loi0iLOloLLL <= 32'hffff_ffff ;
 OoLl0IIIo0IollLoILOLlOIiioIIi0iIo <= 32'hffff_ffff ;
 OIoIi0IlLoooi0iILio0lILiIOL0oLOol <= 32'hffff_ffff ;
 OIlooiLoolLOlLiOLioooILlolIlIlIoi <= 32'hffff_ffff ;
 OiloOOiiooL0o0OIOOiiL0Iii0Lii0LLi <= 32'hffff_ffff ;
 O0O0Il000ILILl0iIOIOOIi00OilLLLoi <= 32'hffff_ffff ;
 OLoi0olioL0OLoILii0iO00IlOOLI00l0 <= 32'hffff_ffff ;
 OOlILI0loI0illoollOiIIOl0iii0oIIi <= 32'hffff_ffff ;
 OiL0iLlILIoiO0lLioo0ololOiILIIoOl <= 32'hffff_ffff ;
 OlllolOIO000iLIo0I0LoLoOLL0IlLl0O <= 32'hffff_ffff ;
 OIIOLlIiiOoLOLLoLOOO0OOoOoOLIOool <= 32'hffff_ffff ;
 OOoLoiLILiiOi0OoO0olOoOoioo0lLoLl <= 32'hffff_ffff ;
 OLiLOi0l0li0loOLOIolIOIIOiLlilolI <= 32'hffff_ffff ;
 OlLIiII0LOiOOo0OoloIILoOIoIOi0O00 <= 32'hffff_ffff ;
 O0OLOILIl0iOLLOoL0LIOIooloLOLo0ii <= 32'hffff_ffff ;
 OLLOi0ioLIIiliILllOIIioOl0OLilili <= 32'hffff_ffff ;
 OLi0IOOoOL00iloIi0i0lLioLiIoioOoo <= 32'hffff_ffff ;
 OIoO0O0OIiIIi00OLLl0olOIOiiIIl0IO <= 32'hffff_ffff ;
 OoIlOlOiL0ollilOlli00LlIOlioLi0l0 <= 32'hffff_ffff ;
 OOllii0LlOLLLoLOIOOiiIO0LlIoooOIL <= 32'hffff_ffff ;
 OoilOILoi0lOli00o0lol0ILilOolil0l <= 32'hffff_ffff ;
 OLOLOILIoOlIiL0iLOooilloILI0OiLlo <= 32'hffff_ffff ;
 O0ooio00O00Ii0l0iill0iLLOLLOOOIIo <= 32'hffff_ffff ;
 OoOOo0iiI0iLoIooI0OIOOiLO0IooOILO <= 32'hffff_ffff ;
 OoIOL0IiLi0i0Loi0llllioOoiIoOLLIo <= 32'hffff_ffff ;
 OliLLl0OlLIiOlIIiLlLlooO0LoiLiooO <= 32'hffff_ffff ;
 OioioLOliOLI0IOlLOolII0L0oi0oIiLO <= 32'hffff_ffff ;
 O0l0LioII0IlliOlIIi0IlI00IoOOoiOo <= 32'hffff_ffff ;
 end
 else if ( O0i00oOl00OoIIOIil0LLOi0looIOIL00 ) begin
 OoloOOilIOLlIlIII0oIL0IOllO0oLi0o <= OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 O0OoOIloiOI0oOil0LlIl0oil0iLOOiLL <= OoloOOilIOLlIlIII0oIL0IOllO0oLi0o ;
 OlLO0OLOOiLioiL0ILLllii0OlIiOOIo0 <= O0OoOIloiOI0oOil0LlIl0oil0iLOOiLL ;
 O0OIlIIlo00lILOO0iOiIILOOI0OI0oOi <= OlLO0OLOOiLioiL0ILLllii0OlIiOOIo0 ;
 O0i0lIILioOLiLOIiIO00loi0iLOloLLL <= O0OIlIIlo00lILOO0iOiIILOOI0OI0oOi ;
 OoLl0IIIo0IollLoILOLlOIiioIIi0iIo <= O0i0lIILioOLiLOIiIO00loi0iLOloLLL ;
 OIoIi0IlLoooi0iILio0lILiIOL0oLOol <= OoLl0IIIo0IollLoILOLlOIiioIIi0iIo ;
 OIlooiLoolLOlLiOLioooILlolIlIlIoi <= OIoIi0IlLoooi0iILio0lILiIOL0oLOol ;
 OiloOOiiooL0o0OIOOiiL0Iii0Lii0LLi <= OIlooiLoolLOlLiOLioooILlolIlIlIoi ;
 O0O0Il000ILILl0iIOIOOIi00OilLLLoi <= OiloOOiiooL0o0OIOOiiL0Iii0Lii0LLi ;
 OLoi0olioL0OLoILii0iO00IlOOLI00l0 <= O0O0Il000ILILl0iIOIOOIi00OilLLLoi ;
 OOlILI0loI0illoollOiIIOl0iii0oIIi <= OLoi0olioL0OLoILii0iO00IlOOLI00l0 ;
 OiL0iLlILIoiO0lLioo0ololOiILIIoOl <= OOlILI0loI0illoollOiIIOl0iii0oIIi ;
 OlllolOIO000iLIo0I0LoLoOLL0IlLl0O <= OiL0iLlILIoiO0lLioo0ololOiILIIoOl ;
 OIIOLlIiiOoLOLLoLOOO0OOoOoOLIOool <= OlllolOIO000iLIo0I0LoLoOLL0IlLl0O ;
 OOoLoiLILiiOi0OoO0olOoOoioo0lLoLl <= OIIOLlIiiOoLOLLoLOOO0OOoOoOLIOool ;
 OLiLOi0l0li0loOLOIolIOIIOiLlilolI <= OOoLoiLILiiOi0OoO0olOoOoioo0lLoLl ;
 OlLIiII0LOiOOo0OoloIILoOIoIOi0O00 <= OLiLOi0l0li0loOLOIolIOIIOiLlilolI ;
 O0OLOILIl0iOLLOoL0LIOIooloLOLo0ii <= OlLIiII0LOiOOo0OoloIILoOIoIOi0O00 ;
 OLLOi0ioLIIiliILllOIIioOl0OLilili <= O0OLOILIl0iOLLOoL0LIOIooloLOLo0ii ;
 OLi0IOOoOL00iloIi0i0lLioLiIoioOoo <= OLLOi0ioLIIiliILllOIIioOl0OLilili ;
 OIoO0O0OIiIIi00OLLl0olOIOiiIIl0IO <= OLi0IOOoOL00iloIi0i0lLioLiIoioOoo ;
 OoIlOlOiL0ollilOlli00LlIOlioLi0l0 <= OIoO0O0OIiIIi00OLLl0olOIOiiIIl0IO ;
 OOllii0LlOLLLoLOIOOiiIO0LlIoooOIL <= OoIlOlOiL0ollilOlli00LlIOlioLi0l0 ;
 OoilOILoi0lOli00o0lol0ILilOolil0l <= OOllii0LlOLLLoLOIOOiiIO0LlIoooOIL ;
 OLOLOILIoOlIiL0iLOooilloILI0OiLlo <= OoilOILoi0lOli00o0lol0ILilOolil0l ;
 O0ooio00O00Ii0l0iill0iLLOLLOOOIIo <= OLOLOILIoOlIiL0iLOooilloILI0OiLlo ;
 OoOOo0iiI0iLoIooI0OIOOiLO0IooOILO <= O0ooio00O00Ii0l0iill0iLLOLLOOOIIo ;
 OoIOL0IiLi0i0Loi0llllioOoiIoOLLIo <= OoOOo0iiI0iLoIooI0OIOOiLO0IooOILO ;
 OliLLl0OlLIiOlIIiLlLlooO0LoiLiooO <= OoIOL0IiLi0i0Loi0llllioOoiIoOLLIo ;
 OioioLOliOLI0IOlLOolII0L0oi0oIiLO <= OliLLl0OlLIiOlIIiLlLlooO0LoiLiooO ;
 O0l0LioII0IlliOlIIi0IlI00IoOOoiOo <= OioioLOliOLI0IOlLOolII0L0oi0oIiLO ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOOLIoiLiLOOLooIoOoioiooIIoliLOlo <= 1'd0 ;
 O0llLOll00OIl0OoLOiOiioIo0O0IolOo <= 1'd0 ;
 OlIiOlLoi0loOiLoLoioiIOIioliiLill <= 1'd0 ;
 OOlL0lLllIOooOI0Ol0L0olliOLO0IlII <= 1'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OOOLIoiLiLOOLooIoOoioiooIIoliLOlo <= 1'd0 ;
 O0llLOll00OIl0OoLOiOiioIo0O0IolOo <= 1'd0 ;
 OlIiOlLoi0loOiLoLoioiIOIioliiLill <= 1'd0 ;
 OOlL0lLllIOooOI0Ol0L0olliOLO0IlII <= 1'd0 ;
 end
 else if ( OllII0i0lILiOLIL0OiIIoLoiIl0IoLoI ) begin
 OOOLIoiLiLOOLooIoOoioiooIIoliLOlo <= ( (OoloOOilIOLlIlIII0oIL0IOllO0oLi0o==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0OoOIloiOI0oOil0LlIl0oil0iLOOiLL==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OlLO0OLOOiLioiL0ILLllii0OlIiOOIo0==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0OIlIIlo00lILOO0iOiIILOOI0OI0oOi==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0i0lIILioOLiLOIiIO00loi0iLOloLLL==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OoLl0IIIo0IollLoILOLlOIiioIIi0iIo==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OIoIi0IlLoooi0iILio0lILiIOL0oLOol==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OIlooiLoolLOlLiOLioooILlolIlIlIoi==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) );
 O0llLOll00OIl0OoLOiOiioIo0O0IolOo <= ( (OiloOOiiooL0o0OIOOiiL0Iii0Lii0LLi==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0O0Il000ILILl0iIOIOOIi00OilLLLoi==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OLoi0olioL0OLoILii0iO00IlOOLI00l0==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OOlILI0loI0illoollOiIIOl0iii0oIIi==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OiL0iLlILIoiO0lLioo0ololOiILIIoOl==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OlllolOIO000iLIo0I0LoLoOLL0IlLl0O==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OIIOLlIiiOoLOLLoLOOO0OOoOoOLIOool==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OOoLoiLILiiOi0OoO0olOoOoioo0lLoLl==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) );
 OlIiOlLoi0loOiLoLoioiIOIioliiLill <= ( (OLiLOi0l0li0loOLOIolIOIIOiLlilolI==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OlLIiII0LOiOOo0OoloIILoOIoIOi0O00==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0OLOILIl0iOLLOoL0LIOIooloLOLo0ii==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OLLOi0ioLIIiliILllOIIioOl0OLilili==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OLi0IOOoOL00iloIi0i0lLioLiIoioOoo==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OIoO0O0OIiIIi00OLLl0olOIOiiIIl0IO==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OoIlOlOiL0ollilOlli00LlIOlioLi0l0==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OOllii0LlOLLLoLOIOOiiIO0LlIoooOIL==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) );
 OOlL0lLllIOooOI0Ol0L0olliOLO0IlII <= ( (OoilOILoi0lOli00o0lol0ILilOolil0l==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OLOLOILIoOlIiL0iLOooilloILI0OiLlo==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0ooio00O00Ii0l0iill0iLLOLLOOOIIo==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OoOOo0iiI0iLoIooI0OIOOiLO0IooOILO==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OoIOL0IiLi0i0Loi0llllioOoiIoOLLIo==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OliLLl0OlLIiOlIIiLlLlooO0LoiLiooO==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (OioioLOliOLI0IOlLOolII0L0oi0oIiLO==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) || (O0l0LioII0IlliOlIIi0IlI00IoOOoiOo==OLo0oiiL0ooIliO0I0illLoILiiIoIoOI) );
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OoILOLi0I0lO0LOI0Illoo0Lo0ilOLLoL <= 1'd0 ;
 end
 else begin
 OoILOLi0I0lO0LOI0Illoo0Lo0ilOLLoL <= OOOLIoiLiLOOLooIoOoioiooIIoliLOlo || O0llLOll00OIl0OoLOiOiioIo0O0IolOo || OlIiOlLoi0loOiLoLoioiIOIioliiLill || OOlL0lLllIOooOI0Ol0L0olliOLO0IlII ;
 end
 end
 wire [31:0] O0ilIlIlLIolLOIIoiooLoiLOiliOOOiO = O0o0loiLIOlLoi0iOIolL0LoOILoilLLl + 1'd1 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0Loo0iiI0OlLOlOIiILOooOOlIoioOli <= 1'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OI00OiLolooiIIiiILoIliO0O0loolIlI) begin
 O0Loo0iiI0OlLOlOIiILOooOOlIoioOli <= 1'd1 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&~OI00OiLolooiIIiiILoIliO0O0loolIlI) begin
 O0Loo0iiI0OlLOlOIiILOooOOlIoioOli <= 1'd0 ;
 end
 else if ( OiliiIIiiIOoIIOOoOo0Oii00ollOOIoO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd12 ) && OliOOOIooO0oILLiLiiilLIlilo0ooL0O ) begin
 if ( (O0ilIlIlLIolLOIIoiooLoiLOiliOOOiO<=OO0liOO0iOOIioool0OoLliiiI0l0ilOo) ) begin
 O0Loo0iiI0OlLOlOIiILOooOOlIoioOli <= 1'd0 ;
 end
 else begin
 O0Loo0iiI0OlLOlOIiILOooOOlIoioOli <= 1'd1 ;
 end
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= 1'd0 ;
 end
 else if (OI0OOlIliLiLli0iiiOOl0lLoOIoLi0Li && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd16) && (OOOi0LIiLLOLIoliiOlolloOli0oLLioi >= (O0oioIoloolL0oiioLILllioiO0oliIOl-1'b1) ) && (Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi==4'd0) && (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) ) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= OliOOOIooO0oILLiLiiilLIlilo0ooL0O && ( OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 || OI00liOIoliolOollOLoioOLooloiloI0 ) && ~OoILOLi0I0lO0LOI0Illoo0Lo0ilOLLoL ;
 end
 else if (OOIIIOLL0O000ioLliOIoOii0LiI0lOoo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oi0lIlIOooiiiI0I00Ol0ioiiL0liiOIi) && (OliiLIIliIO0OIloloLiiI0ilOILLILOI>=OILLIiOoiIOiIil0OLOLLiIIllIlOLilI) ) begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= OliOOOIooO0oILLiLiiilLIlilo0ooL0O && ( OLOlLL0i0OIOoLIOIlLiIiLlOOllOO0l0 || OI00liOIoliolOollOLoioOLooloiloI0 ) && ~OoILOLi0I0lO0LOI0Illoo0Lo0ilOLLoL;
 end
 else begin
 O0i00oOl00OoIIOIil0LLOi0looIOIL00 <= 1'd0 ;
 end
 end
 reg [47:0] OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl <= 48'd0 ;
 OOOll0oL0OOLoi0lIioOo0liiLILLoiiL <= 1'd0 ;
 end
 else if ( OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) begin
 OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl <= 48'd0 ;
 OOOll0oL0OOLoi0lIioOo0liiLILLoiiL <= 1'd0 ;
 end
 else if ( O0i00oOl00OoIIOIil0LLOi0looIOIL00 ) begin
 OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl <= 48'd0 ;
 OOOll0oL0OOLoi0lIioOo0liiLILLoiiL <= 1'd0 ;
 end
 else if ( (OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl>({OoIolioOL0iLLOLloI00iIILLiiL0Ooil,16'hffff})) && OiiLOILl0iLi0L0ilIIoooLLIoliIIIlO ) begin
 OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl <= 48'd0 ;
 OOOll0oL0OOLoi0lIioOo0liiLILLoiiL <= 1'd1 ;
 /* synthesis translate_off */ $display("%m Warning OOOll0oL0OOLoi0lIioOo0liiLILLoiiL !!!!! \n " );
 /* synthesis translate_on */ end
 else begin
 OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl <= (OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl==48'hffff_ffff_ffff) ? OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl : OiLOOO0iiLiiOLIoLIIOIi0LoOO0I0LIl + 64'd1 ;
 OOOll0oL0OOLoi0lIioOo0liiLILLoiiL <= 1'd0 ;
 end
 end
 OoLiL0iillLiLlLlO0loIIoLl0l0l0LoI sq_fir_cut_out ( .OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ( OOllOo00o0IlooI0l0io0O00l0OIoiILO ), .OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ( OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ), .OI00OiLolooiIIiiILoIliO0O0loolIlI ( OOL0o0i0Llo0IiiLlO00oliOILLI00Ool ), .O0Loo0iiI0OlLOlOIiILOooOOlIoioOli (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ), .O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo (O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ) , .OILIloOoilLIL00IIOoOilLOO0L0iiIOO (OILIloOoilLIL00IIOoOilLOO0L0iiIOO), .O0oLLi0Ill00l0lioiLioiooIllloIiIl (O0oLLi0Ill00l0lioiLioiooIllloIiIl), .OilOIloOO0LiLoIL0IIILoIi0Loilll0I (OilOIloOO0LiLoIL0IIILoIi0Loilll0I ), .Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 (Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ), .OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O (OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ), .OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO (OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ), .OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 (OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ), .OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ( OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ) , .OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ( OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ) , .OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ( OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ) , .OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ( OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ) , .OiooiLLioLLL0lII00ol0oIOllLlOiLlL ( OiooiLLioLLL0lII00ol0oIOllLlOiLlL ) , .OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ( OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ) , .O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ( O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ) , .Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ( Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ) , .O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ( O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ) , .OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ( OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ) , .OilLIO0lI0LO0LolOOilILl0oiIlolOlo ( OilLIO0lI0LO0LolOOilILl0oiIlolOlo ) , .OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ( OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ) , .OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ( OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ) , .OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ( OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ) , .OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ( OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ) , .OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ( OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ) , .OIoliiOo0i000ooilOOLOiil0LlLiOoLo ( OIoliiOo0i000ooilOOLOiil0LlLiOoLo ) , .Oo00OlooOo0io0OoIloiioLiOlL0llio0 ( Oo00OlooOo0io0OoIloiioLiOlL0llio0 ) , .OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ( OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ) , .OOoOoILioOoIlIoLliOLOOi0io0IlLolo ( OOoOoILioOoIlIoLliOLOOi0io0IlLolo ) , .OiLllooo0Li0lioiolLi0ILIoLOliil0I ( OiLllooo0Li0lioiolLi0ILIoLOliil0I ) , .OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ( OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ) , .OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ( OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ) , .OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ( OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ) , .OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ( OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ) , .OLL0OiLILloil0IoOlLIIloLIiIlllLil ( OLL0OiLILloil0IoOlLIIloLIiIlllLil ) , .OILI0LLillilOlllLil0ioLoIiliOoLLo ( OILI0LLillilOlllLil0ioLoIiliOoLLo ) , .OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ( OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ) , .OoIloII0oLiOLOLIllOL0iOoooOliOIii ( OoIloII0oLiOLOLIllOL0iOoooOliOIii ) , .Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ( Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ) , .OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ( OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ) , .O0oill0llILOilo0i0LIoOLIoolL0Il0o (O0oill0llILOilo0i0LIoOLIoolL0Il0o ), .OlliILlLOilOl0LO0O0OilooiIIiOi0Ll (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ), .OiL0LolLLIOlliloII00llOil0oIlOiIo (OiL0LolLLIOlliloII00llOil0oIlOiIo ), .O0llIOIliLOO0iiOoO0OO0lIOloLoII0I (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I), .OOLoL0looIOoioIoOooIoLIiIiLiLoiOl (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ), .OIoIooIolOilIOlooOlOIIOoilLioOIIO (OIoIooIolOilIOlooOlOIIOoilLioOIIO ), .Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] ), .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ), .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl ), .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 (OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ), .O0lOIlooLi0lilOllLlilIo00iOLiOLLo (O0lOIlooLi0lilOllLlilIo00iOLiOLLo ), .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo ), .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) );
 OLiIILolLli0LiLoOOo0lIlOiOoO0lioL OLiIILolLli0LiLoOOo0lIlOiOoO0lioL ( .OOLIiil0IlIllLollIl0LIilliOI0iolo (OOLIiil0IlIllLollIl0LIilliOI0iolo ) , .O0il0IO0olIoLiOIL0000lo0OoliIL0Ll (O0il0IO0olIoLiOIL0000lo0OoliIL0Ll ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI (OOLOoolOi0LIo0olO0loLllIlllIiiIiI ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI (OOOLiLOilooIi0Iio00ilILoLIILOoOoI ) , .OLLOooI0ILL00ILloiliILLLiioooLliI (OLLOooI0ILL00ILloiliILLLiioooLliI ) , .OL0O0IIio0loL0L0Il0li0i00lliIoOOI (OL0O0IIio0loL0L0Il0li0i00lliIoOOI ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI (OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ) , .Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ) , .O0lOIlooLi0lilOllLlilIo00iOLiOLLo (O0lOIlooLi0lilOllLlilIo00iOLiOLLo ) , .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ) , .Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl (Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ) , .O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI (O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ) , .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) );
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIloLiiOL00oilLo0iiILoOOll0lIlIlO <= 32'd0 ;
 end
 else begin
 OIloLiiOL00oilLo0iiILoOOll0lIlIlO <= {24'd0,3'd0 , (OiiLOILl0iLi0L0ilIIoooLLIoliIIIlO&&~Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII) , OlIl0ooIoiLlO0lII0loOOi0IoIILloOO||OiLoLOLiLooLLi0loLlLiooo0LliOiIoL , O0il0IO0olIoLiOIL0000lo0OoliIL0Ll , OOooLlloIiioOOO0LLILl0liiillLILol , O0IIOOO0LOOiLiiOill00LllllIOIILo0 } ;
 end
 end
 endmodule
 module OILLilL0iiliiLLO0IL0LiOoLILlOL0iO ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L , OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl , OoIolioOL0iLLOLloI00iIILLiiL0Ooil , OOLIiil0IlIllLollIl0LIilliOI0iolo, OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI , OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 , OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI, , OilOOo00lLiOOoiO0ii0oo0oOliOollii, , OLll00OOliOil0O0iLlIooLOLooIIlI0o, O0o0loiLIOlLoi0iOIolL0LoOILoilLLl, OO0liOO0iOOIioool0OoLliiiI0l0ilOo, OiIOLi00lOILlOOL0oLLloL0io0LoIoOL, OolIOLOooiLLIllI0LOLIolllLoilolIl , O0IOooLliOlIllOliILoolIIoIiO0Ilol , OLo0oiiL0ooIliO0I0illLoILiiIoIoOI , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 , OoiloolOiOIoIOolLiOl0OlOiOli0oOOl , OillLliLoolOIiiiILoOILOIloo000iLI , OlLOLoI0iIOLloliOllILlOoIiioOli0L , OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI , OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII , OOLOoolOi0LIo0olO0loLllIlllIiiIiI , OOOLiLOilooIi0Iio00ilILoLIILOoOoI , OLLOooI0ILL00ILloiliILLLiioooLliI , OILoli0OIOIIOI0OiliOo0i0OLoliOOiI , O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI , OL0O0IIio0loL0L0Il0li0i00lliIoOOI , OilOOioILlOIIOL0iioIOIi0oloooOoLl , OI00OiLolooiIIiiILoIliO0O0loolIlI , OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo , OIloLiiOL00oilLo0iiILoOOll0lIlIlO , OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O , OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI , OIIOLLOIlOlLoi0oiOioLilOiioiiliLO , OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi, OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 , Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL, OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI );
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input [3:0] Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L ;
 input [3:0] OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl ;
 input [31:0] OoIolioOL0iLLOLloI00iIILLiiL0Ooil ;
 output [4:0] OOLIiil0IlIllLollIl0LIilliOI0iolo;
 output [31:0] OLll00OOliOil0O0iLlIooLOLooIIlI0o;
 output [31:0] O0o0loiLIOlLoi0iOIolL0LoOILoilLLl;
 output [31:0] OO0liOO0iOOIioool0OoLliiiI0l0ilOo;
 output OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 input [ 15: 0] OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ;
 output [31:0] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 input [15:0] OoiloolOiOIoIOolLiOl0OlOiOli0oOOl ;
 input [15:0] OillLliLoolOIiiiILoOILOIloo000iLI ;
 input [15:0] OlLOLoI0iIOLloliOllILlOoIiioOli0L ;
 input OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ;
 input [ 3: 0] OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 input OOLOoolOi0LIo0olO0loLllIlllIiiIiI ;
 input OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 input [ 63: 0] OLLOooI0ILL00ILloiliILLLiioooLliI ;
 input [ 2: 0] OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 input [ 15: 0] O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ;
 output OL0O0IIio0loL0L0Il0li0i00lliIoOOI ;
 input [ 15: 0] OilOOioILlOIIOL0iioIOIi0oloooOoLl ;
 input [31:0] OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 input [31:0] OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ;
 output [31:0] OIloLiiOL00oilLo0iiILoOOll0lIlIlO ;
 output [31:0] OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ;
 output [31:0] OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ;
 input [ 15: 0] OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ;
 output OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi;
 output [255:0] OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 ;
 output Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL;
 input OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI;
 wire [31:0] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 wire [31:0] OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ;
 wire [31:0] O0I0oI0I000LllOOI0L0lOlIl000LIioO ;
 wire Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ;
 wire O0oill0llILOilo0i0LIoOLIoolL0Il0o ;
 wire OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ;
 wire OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ;
 wire OIoIooIolOilIOlooOlOIIOoilLioOIIO ;
 wire OiL0LolLLIOlliloII00llOil0oIlOiIo ;
 wire O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ;
 wire OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL ;
 wire [31:0] OilOIloOO0LiLoIL0IIILoIi0Loilll0I ;
 wire [31:0] Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ;
 wire [31:0] OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ;
 wire [63:0] OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ;
 wire [ 2:0] OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ;
 wire [ 2:0] OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ;
 wire [ 2:0] OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ;
 wire [ 2:0] OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ;
 wire [ 2:0] OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ;
 wire [ 2:0] OiooiLLioLLL0lII00ol0oIOllLlOiLlL ;
 wire [ 2:0] OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ;
 wire [ 2:0] O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ;
 wire [ 2:0] Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ;
 wire [ 2:0] O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ;
 wire [ 2:0] OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ;
 wire [ 2:0] OilLIO0lI0LO0LolOOilILl0oiIlolOlo ;
 wire [ 2:0] OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ;
 wire [ 2:0] OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ;
 wire [ 2:0] OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ;
 wire [ 2:0] OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ;
 wire [ 2:0] OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ;
 wire [ 2:0] OIoliiOo0i000ooilOOLOiil0LlLiOoLo ;
 wire [ 2:0] Oo00OlooOo0io0OoIloiioLiOlL0llio0 ;
 wire [ 2:0] OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ;
 wire [ 2:0] OOoOoILioOoIlIoLliOLOOi0io0IlLolo ;
 wire [ 2:0] OiLllooo0Li0lioiolLi0ILIoLOliil0I ;
 wire [ 2:0] OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ;
 wire [ 2:0] OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ;
 wire [ 2:0] OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ;
 wire [ 2:0] OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ;
 wire [ 2:0] OLL0OiLILloil0IoOlLIIloLIiIlllLil ;
 wire [ 2:0] OILI0LLillilOlllLil0ioLoIiliOoLLo ;
 wire [ 2:0] OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ;
 wire [ 2:0] OoIloII0oLiOLOLIllOL0iOoooOliOIii ;
 wire [ 2:0] Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ;
 wire [ 2:0] OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ;
 wire [31:0] O0o0loiLIOlLoi0iOIolL0LoOILoilLLl = 32'd0 ;
 wire [31:0] OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 wire OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 wire [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 wire [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 wire [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 wire [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 wire [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 wire [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 wire [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 wire [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 wire [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 wire [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 wire [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 wire [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 wire [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 wire [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 wire [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 wire [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 wire O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 wire [ 23: 0] OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ;
 wire [ 23: 0] OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ;
 wire [ 23: 0] O0oLiillllLOiLilOoI000iOLoiL0L0LO ;
 wire [ 23: 0] Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ;
 wire [ 23: 0] OoooIiooOl0i0oliO0lio0IOo0iIILLLi ;
 wire [ 23: 0] OLlLoL0lO0oOIOolIIoiILIO0oOilooll ;
 wire [ 23: 0] OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ;
 wire [ 23: 0] Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ;
 wire [ 23: 0] Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ;
 wire [ 23: 0] OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ;
 wire [ 23: 0] Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ;
 wire [ 23: 0] OLi0ooOo0OlIllLOILllLL00lL00Liii0 ;
 wire [ 23: 0] OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ;
 wire [ 23: 0] OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ;
 wire [ 23: 0] OOIlIio0iILll00lliIIioiIiOLlLLi00 ;
 wire [ 23: 0] OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ;
 wire [ 23: 0] OLio000LoL0lOol0oIiLlILLIlOLLOIlO ;
 wire [ 23: 0] OoiiooOo00OI0O0loiolLOLioIOiI0LoI ;
 wire [ 23: 0] Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ;
 wire [ 23: 0] OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ;
 wire [ 23: 0] OIO0IioIOoIOIll0LOIlOOILoILoiilli ;
 wire [ 23: 0] OLoOLiILLLiIilOolo0Lil0iLLOOLILII ;
 wire [ 23: 0] OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ;
 wire [ 23: 0] OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ;
 wire [ 23: 0] OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ;
 wire [ 23: 0] OlIli0IolOiL0LoliLloo0olllliIiO0O ;
 wire [ 23: 0] OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ;
 wire [ 23: 0] Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ;
 wire [ 23: 0] OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ;
 wire [ 23: 0] OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ;
 wire [ 23: 0] OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ;
 wire [ 23: 0] O0lolLi0olIioIiIooOLLLlioIooLIill ;
 wire [ 7: 0] OoolLolOioLILoOIII00LIOli00LIlloi ;
 wire [ 7: 0] OOIolooo0Oi00io00lIiiOiiLIliliOio ;
 wire [ 7: 0] OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ;
 wire [ 7: 0] OOoL0lOOloLLOLOILLLOolliIll0oOOoO ;
 wire [ 7: 0] OoOlILlliliiOI0OLLoOOl0000iIo0IIo ;
 wire [ 7: 0] O0iI0Lil0liLOLiILLOoilII0LII0iolO ;
 wire [ 7: 0] O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ;
 wire [ 7: 0] O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ;
 wire [ 7: 0] O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ;
 wire [ 7: 0] OIO0IIi0OIooOiLOIII0lLolililiOIll ;
 wire [ 7: 0] OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ;
 wire [ 7: 0] OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ;
 wire [ 7: 0] OO0OOoLL0O0OOOllioILi0liilLLloiLO ;
 wire [ 7: 0] OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ;
 wire [ 7: 0] OlIollIiLi0IlLiolloLOOL000Oo0l0II ;
 wire [ 7: 0] O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ;
 wire [ 7: 0] OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ;
 wire [ 7: 0] OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ;
 wire [ 7: 0] OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ;
 wire [ 7: 0] O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ;
 wire [ 7: 0] Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ;
 wire [ 7: 0] O00liliooOOoiI0OlOOIIlO0o0IiOOolL ;
 wire [ 7: 0] O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ;
 wire [ 7: 0] Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ;
 wire [ 7: 0] OlLIiOlioIILOllO00lLiI0LiIlOloIiI ;
 wire [ 7: 0] OO00il0IO0lLoiilIo0ioiOiOOlLloioL ;
 wire [ 7: 0] OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ;
 wire [ 7: 0] O0oIiILIIO0LOOil00IlIoLiIilO00ooI ;
 wire [ 7: 0] OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ;
 wire [ 7: 0] OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ;
 wire [ 7: 0] OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ;
 wire [ 7: 0] OolLO0OOloooOIOiiOilL0IiILL0iol0I ;
 wire [ 31: 0] OOOooLlOLO0iOOOLi00oIiloILlooOLIO ;
 wire [ 31: 0] OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ;
 wire [ 31: 0] Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ;
 wire [ 31: 0] OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ;
 wire [ 31: 0] OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ;
 wire [ 31: 0] OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ;
 wire [ 31: 0] OoLLliL00LLoooll00ooiLolOliOO0lLI ;
 wire [ 31: 0] O0li0llLIi0oIo0IilLLooLILolLIOOoo ;
 wire [ 31: 0] OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ;
 wire [ 31: 0] OioilLoll0OiiOooiLiIOiL0LiilILII0 ;
 wire [ 31: 0] Ol0OLoIiI0OloLIlillLOloLioIIL0III ;
 wire [ 31: 0] Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ;
 wire [ 31: 0] OlLlliliOioioOIoiLOIOiOoiiioIOLOO ;
 wire [ 31: 0] OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ;
 wire [ 31: 0] OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ;
 wire [ 31: 0] OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ;
 wire [ 31: 0] OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ;
 wire [ 31: 0] O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ;
 wire [ 31: 0] O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ;
 wire [ 31: 0] OO0llOooLooLoi0l0oIOOoilOolIoLLOo ;
 wire [ 31: 0] OLl0oiiIOL0ol00LIoo0IoolIollol0ii ;
 wire [ 31: 0] OILLl0iillioLoOiiIiL0iliIOiO0oiio ;
 wire [ 31: 0] OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ;
 wire [ 31: 0] OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ;
 wire [ 31: 0] OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ;
 wire [ 31: 0] OLoLOlol00olO0oo0LLlolI0OiLo0llLI ;
 wire [ 31: 0] OLolOilolLoloilIloOOiioIloiI0L0Lo ;
 wire [ 31: 0] OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ;
 wire [ 31: 0] OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ;
 wire [ 31: 0] OLololIl0LoiLooLIloiooLli0LOOLLli ;
 wire [ 31: 0] OIllOIIOiOol000OoLIL0lLl0L00iIIIL ;
 wire [ 31: 0] OL0looio0Loioi0ill0olOo0o00ioOOII ;
 wire [ 7: 0] OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ;
 wire [ 7: 0] O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ;
 wire [ 7: 0] OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ;
 wire [ 7: 0] OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ;
 wire [ 7: 0] O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ;
 wire [ 7: 0] OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ;
 wire [ 7: 0] OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ;
 wire [ 7: 0] OioIOIo0IllIo0OILLlli0LOOl00lioII ;
 wire [ 7: 0] O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ;
 wire [ 7: 0] OLoli0Li0i0oO0olOOilIliIio0LOoIIO ;
 wire [ 7: 0] OiILooool0OiolIOIIlO0LiOliIiIL0Ii ;
 wire [ 7: 0] OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ;
 wire [ 7: 0] OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ;
 wire [ 7: 0] O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ;
 wire [ 7: 0] OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ;
 wire [ 7: 0] OOoLol0oioL0looOlO0io0oIillil0iI0 ;
 wire [ 7: 0] OILIi00LOILOoLIiLloLiLIolliOoooIo ;
 wire [ 7: 0] OIi0liIIIoiOooLllLO0O0IoLLllIOlli ;
 wire [ 7: 0] O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ;
 wire [ 7: 0] OOIIlilOoOlIolLlILLioil0LL0oLlloo ;
 wire [ 7: 0] OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ;
 wire [ 7: 0] OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ;
 wire [ 7: 0] OOiOiIiiilililLoLlIOoIoiILilLoooI ;
 wire [ 7: 0] OO0O00OIoioOIOLi0IlILI0OlilooOIOo ;
 wire [ 7: 0] OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ;
 wire [ 7: 0] OlIiO0llI0O0Li00OLIILiOLi00OiLioL ;
 wire [ 7: 0] O0lIlL0lLL00000ioioloooIoiiiioi00 ;
 wire [ 7: 0] OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ;
 wire [ 7: 0] OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ;
 wire [ 7: 0] OILllI0lillIoilOIoooOll0LII00I0l0 ;
 wire [ 7: 0] OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ;
 wire [ 7: 0] Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ;
 wire [ 31: 0] OioLioLloIiilLLoOlIoiLIO0IOoiLoll ;
 wire [ 31: 0] OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ;
 wire [ 31: 0] OI0ioOlloiIio0oiOloi0lioiILoollLl ;
 wire [ 31: 0] O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ;
 wire [ 31: 0] OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ;
 wire [ 31: 0] O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ;
 wire [ 31: 0] O00loOoIIlII0OOo0lio00iOOOolLiIiO ;
 wire [ 31: 0] OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ;
 wire [ 31: 0] O0il0OIIioo0IoL0OI0llOiLiLioill0i ;
 wire [ 31: 0] OLLOoOIo0oiL0IOOO0lill0iloILllIOO ;
 wire [ 31: 0] OlLiiOLII0io0OLOOiIiiO0IIililoolo ;
 wire [ 31: 0] Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ;
 wire [ 31: 0] OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ;
 wire [ 31: 0] OoLiLLooILIo0iol0OIoliLi0iiioiIlI ;
 wire [ 31: 0] OiiooiLLOL0iiO0oILoOlLoololiIIo0o ;
 wire [ 31: 0] OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ;
 wire [ 31: 0] OioilI0Oo0oOil0lIioiILIOLLLOLLioO ;
 wire [ 31: 0] OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ;
 wire [ 31: 0] O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ;
 wire [ 31: 0] OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ;
 wire [ 31: 0] OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ;
 wire [ 31: 0] O0I0LooLLiIO0illo0IliLLoioL0LlOLl ;
 wire [ 31: 0] OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ;
 wire [ 31: 0] OlLo00LioOiOOOoliolIoLI0olOOlLoOI ;
 wire [ 31: 0] OliiLi0oooOIo0L0lLoil0ooooi00I0ol ;
 wire [ 31: 0] OoL0LLOIlII0oLlloILillo0IOilOi0Il ;
 wire [ 31: 0] Oioo00O0OIloLlOil00lLiI0oIOOOoIio ;
 wire [ 31: 0] OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ;
 wire [ 31: 0] O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ;
 wire [ 31: 0] OLiILL00lIlOliLloi0OOl00LlIl0Loli ;
 wire [ 31: 0] OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ;
 wire [ 31: 0] Ol0LioliiiiOil0liLiOiolioOo0oioii ;
 wire [175: 0] Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ;
 wire [175: 0] OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ;
 wire [175: 0] OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ;
 wire [175: 0] OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ;
 wire [175: 0] OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ;
 wire [175: 0] OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ;
 wire [175: 0] OiiOIoolI0LioIo0IlL0lOllILIOOiIio ;
 wire [175: 0] OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ;
 wire [175: 0] O0lioOi00lO0IL00IoLLILolIlli00LiI ;
 wire [175: 0] OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ;
 wire [175: 0] OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ;
 wire [175: 0] Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ;
 wire [175: 0] OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ;
 wire [175: 0] OI0ool0i0ollOOoloL00L0LlLIO0LIliI ;
 wire [175: 0] OL0Lio0lIililolilllOL0Li0lIi0I0LI ;
 wire [175: 0] OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ;
 wire [175: 0] OI0L0iIOilOi0LlILL0l0liiiil0lOIii ;
 wire [175: 0] OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ;
 wire [175: 0] OooOIi00Ii0liOollOoLioI0OiLiLiO0O ;
 wire [175: 0] OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ;
 wire [175: 0] OiILIII00lOolOiililIOiIIloo0OlLlo ;
 wire [175: 0] OiioOooilOllI0oOoolilo0OLIlioo0II ;
 wire [175: 0] OIiolOOI00iliL0LolLOOOLOliiIlLlII ;
 wire [175: 0] OLOL0OioiLOLoli0LOL00OOiO0iiOooll ;
 wire [175: 0] O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ;
 wire [175: 0] OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ;
 wire [175: 0] O0oL00LOlilLooOoiil0oLL0iIillLlLL ;
 wire [175: 0] Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ;
 wire [175: 0] OIOio00oLLL0o00LO00LLoI0LlL0OILlO ;
 wire [175: 0] OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ;
 wire [175: 0] OlLiolooLilLlLiil0l0iiO0IOILool00 ;
 wire [175: 0] Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ;
 wire [ 71: 0] OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ;
 wire [ 71: 0] Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ;
 wire [ 71: 0] OlIloooO00OIL0L0iIili0iOOoiLI0oiI ;
 wire [ 71: 0] O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ;
 wire [ 71: 0] OLolLol0lLIIlIillI000oIlilLLloOii ;
 wire [ 71: 0] OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ;
 wire [ 71: 0] OoIooolIllLIIolLII0IiLLiiOlOOIIOO ;
 wire [ 71: 0] Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ;
 wire [ 71: 0] OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ;
 wire [ 71: 0] OIILOOOOIOl00OoIollioiiliIilolLLl ;
 wire [ 71: 0] OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ;
 wire [ 71: 0] OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ;
 wire [ 71: 0] OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ;
 wire [ 71: 0] Oo0loliLllliloIiliOi0lILloLI0ILlO ;
 wire [ 71: 0] O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ;
 wire [ 71: 0] O0oilLoOiOiLLi0Li0lLOIooIiliILlii ;
 wire [ 71: 0] OlIIioIIlILoli0oIiIl0l0IlOlloooll ;
 wire [ 71: 0] OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ;
 wire [ 71: 0] OioolLOlII0IlolOIiLOliilL0oiiOoIo ;
 wire [ 71: 0] OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ;
 wire [ 71: 0] OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ;
 wire [ 71: 0] OIolOIIiLIloloOL0iIIO0il0li00ilOo ;
 wire [ 71: 0] O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ;
 wire [ 71: 0] OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ;
 wire [ 71: 0] OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ;
 wire [ 71: 0] OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ;
 wire [ 71: 0] OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ;
 wire [ 71: 0] OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ;
 wire [ 71: 0] OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ;
 wire [ 71: 0] OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ;
 wire [ 71: 0] OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ;
 wire [ 71: 0] OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ;
 wire [ 31: 0] OIiO0OLioLiIOIIiLoiLooI00I0olI00O ;
 wire [ 31: 0] O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ;
 wire [ 31: 0] OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ;
 wire [ 31: 0] O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ;
 wire [ 31: 0] OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ;
 wire [ 31: 0] OLLloO00IliLiLLlLloLloO0liOoIIOOI ;
 wire [ 31: 0] OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ;
 wire [ 31: 0] OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ;
 wire [ 31: 0] OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ;
 wire [ 31: 0] OiooooLLoI0OLilIIil0ilooLo0OIloLl ;
 wire [ 31: 0] OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ;
 wire [ 31: 0] OOOLilOolI0LILLIoloIiO00OiIiLiiIo ;
 wire [ 31: 0] OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ;
 wire [ 31: 0] Ooi0OL0i0IioliooLiI00OoiL00looOIL ;
 wire [ 31: 0] OolL0oo00LOo0LOoLiILllLo0loOoIiii ;
 wire [ 31: 0] O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ;
 wire [ 31: 0] O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ;
 wire [ 31: 0] OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ;
 wire [ 31: 0] OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ;
 wire [ 31: 0] OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ;
 wire [ 31: 0] OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ;
 wire [ 31: 0] OlOllIloiIIIIloliooOo0LoIil0o0oii ;
 wire [ 31: 0] O0OoiooiIOLOllil0OLoLOlllL000LII0 ;
 wire [ 31: 0] O0oiOOLLiiillOliOOOllO0iO000OOoLI ;
 wire [ 31: 0] OlIIloOL0iLIOLlOlLILlloiioloooILi ;
 wire [ 31: 0] OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ;
 wire [ 31: 0] OOILlooOIliLloiliIOi00LIlLIoli000 ;
 wire [ 31: 0] OiIL00IOiOiiI00oiio0lLOlooIiLiOio ;
 wire [ 31: 0] O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ;
 wire [ 31: 0] OilIl00OOIloIli0LIIii00LIIlILiL0L ;
 wire [ 31: 0] OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ;
 wire [ 31: 0] OO0oIOllioLiLlLLlii0ilL0OlIliIilO ;
 wire [ 63: 0] OOOo0I0LlloiIl0i0il0OLiOlooOOolil ;
 wire [ 63: 0] OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ;
 wire [ 63: 0] OolIilIL0iooOLllOLloloOIlLIiOoLo0 ;
 wire [ 63: 0] OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ;
 wire [ 63: 0] OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ;
 wire [ 63: 0] OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ;
 wire [ 63: 0] OLL0i00LllLlio0oLOLooIL0ilLLllil0 ;
 wire [ 63: 0] OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ;
 wire [ 63: 0] OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ;
 wire [ 63: 0] O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ;
 wire [ 63: 0] OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ;
 wire [ 63: 0] OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ;
 wire [ 63: 0] OliliILl0LLiioool00L00LoLLILio0lO ;
 wire [ 63: 0] OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ;
 wire [ 63: 0] OIOIOlilIolIlLOLlLlll0IiOIiILiOol ;
 wire [ 63: 0] OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ;
 wire [ 63: 0] OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ;
 wire [ 63: 0] OI0OLOILiOlOoolLIilooolollLLo0OOO ;
 wire [ 63: 0] OoII0il0iLlL00iIo0I0OoloiiilLOLIo ;
 wire [ 63: 0] Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ;
 wire [ 63: 0] OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ;
 wire [ 63: 0] OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ;
 wire [ 63: 0] Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ;
 wire [ 63: 0] OIliOOilOillIo00oiOOLIOiLolIIooOl ;
 wire [ 63: 0] OolOOLl0OlII0OiiloIloOO00IllliiLO ;
 wire [ 63: 0] O0o0OillO0LllooIiILLoilol0lii0liL ;
 wire [ 63: 0] OLOlILilLoI0liOiooL00OOlo0i0LiiiI ;
 wire [ 63: 0] OOIIilloi0OiOoo0iI0LI0LI00oILiLio ;
 wire [ 63: 0] OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ;
 wire [ 63: 0] OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ;
 wire [ 63: 0] OIoolOll00LlI00l0oIOLLIOI0I0LIILo ;
 wire [ 63: 0] OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ;
 wire [ 31: 0] OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ;
 wire [ 31: 0] OoI00LooIIlIIlIOOLIoloilI0OoIILLi ;
 wire [ 31: 0] OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ;
 wire [ 31: 0] OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ;
 wire [ 31: 0] OO0O0oOlliIoIOlooIO0lOLolIilLllIO ;
 wire [ 31: 0] OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ;
 wire [ 31: 0] OOiOiOIIoOii0oOLlI0OliIi0liioLLII ;
 wire [ 31: 0] O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ;
 wire [ 31: 0] OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ;
 wire [ 31: 0] OiLiiLILIoLilioiLolliOl0LI00LLil0 ;
 wire [ 31: 0] OLlolloLliiLO0IlIlLo0lIiiloL00OOL ;
 wire [ 31: 0] OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ;
 wire [ 31: 0] OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ;
 wire [ 31: 0] OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ;
 wire [ 31: 0] OiloLLIlO00Il0oo0io0Iilliiil0OolO ;
 wire [ 31: 0] OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ;
 wire [ 31: 0] OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ;
 wire [ 31: 0] O0Il0L0lLloiIiliL0000o0oIOLLILool ;
 wire [ 31: 0] OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ;
 wire [ 31: 0] OOoooLL0l0llOLI0o0oO00LIoLO00LILO ;
 wire [ 31: 0] OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ;
 wire [ 31: 0] OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ;
 wire [ 31: 0] OOl0i0OIIooLiI0IioL0LLILIloOlOllL ;
 wire [ 31: 0] OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ;
 wire [ 31: 0] O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ;
 wire [ 31: 0] OIO0L0iO0iLllOLILO0IoLliLolI00lLI ;
 wire [ 31: 0] O0oOLILIoIlLOIIollLOoL00o0O00OiOo ;
 wire [ 31: 0] Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ;
 wire [ 31: 0] OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ;
 wire [ 31: 0] OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ;
 wire [ 31: 0] OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ;
 wire [ 31: 0] OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ;
 wire [ 63: 0] OLlOlii00IoIl00oIioIiIool0lLiOoLo ;
 wire [ 63: 0] OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ;
 wire [ 63: 0] OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ;
 wire [ 63: 0] Ol000OloII0LlIII00IIOIlOiioOo0Iii ;
 wire [ 63: 0] O00I0iOoILll0oILl0ILloii0LIIOOiIO ;
 wire [ 63: 0] OO00IIiOlOioiOLIiIloilLII0lLL0OOi ;
 wire [ 63: 0] OlOl0iOIioolOiill0OLOloOoLiIlllol ;
 wire [ 63: 0] OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ;
 wire [ 63: 0] OioOlIooLl0IL0LiioIlILIolO0o0ii0l ;
 wire [ 63: 0] Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ;
 wire [ 63: 0] OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ;
 wire [ 63: 0] OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ;
 wire [ 63: 0] OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ;
 wire [ 63: 0] OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ;
 wire [ 63: 0] O0oOL0illOloooo0ioIiOLOooLILllLl0 ;
 wire [ 63: 0] OLiILioillIololIOILoOLlI0LILLliIL ;
 wire [ 63: 0] Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ;
 wire [ 63: 0] OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ;
 wire [ 63: 0] Oi0Liloll0L00OiL0iLli0LO00iloIoLi ;
 wire [ 63: 0] OoilLIlliloO0LoOL00IILioiolLIloi0 ;
 wire [ 63: 0] OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ;
 wire [ 63: 0] OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ;
 wire [ 63: 0] OOOlLolILloIii0oollOil0lI0OOoOoo0 ;
 wire [ 63: 0] OIlOIiiliIlIOIlilliilOl0iILIOOOLO ;
 wire [ 63: 0] OIliolloLooOi0OolOOi0ILOlIliLi0o0 ;
 wire [ 63: 0] OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ;
 wire [ 63: 0] O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ;
 wire [ 63: 0] OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ;
 wire [ 63: 0] O0illollo0oliIl0OolOoIlIILL0OIioO ;
 wire [ 63: 0] OoOoIOoI0LILoIlIliLIioOooOOOIOoli ;
 wire [ 63: 0] OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ;
 wire [ 63: 0] OLOllOoI0IolOloolLolO0lIiolLiIILi ;
 wire [ 63: 0] OIollo0oLlLiI0IILOO00illIILLIoo0o ;
 wire [ 63: 0] O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ;
 wire [ 63: 0] O0lIOiilLOiIOollILlioiiOOiiLOO00i ;
 wire [ 63: 0] OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ;
 wire [ 63: 0] OlolloloolOo0o0LLLIl00Li0iiLl00ol ;
 wire [ 63: 0] OOLIlLlLIloIOoooilolooLloIi0OiiIi ;
 wire [ 63: 0] OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ;
 wire [ 63: 0] OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ;
 wire [ 63: 0] OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ;
 wire [ 63: 0] Oloo0IIooolliliLOLoLoL0oI0LOliLlL ;
 wire [ 63: 0] O00oIiiOLOoilolOol0OIIOII00lllOIo ;
 wire [ 63: 0] OlLi0LOI0LoLioI0loilIlo00iliILIoi ;
 wire [ 63: 0] OLioIOLOILilililoO0ililOi0oiIoo0o ;
 wire [ 63: 0] OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ;
 wire [ 63: 0] Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ;
 wire [ 63: 0] OoOOillllIiloIOIILO0lL0LIl0iOlIII ;
 wire [ 63: 0] OIOO0oiiIiiOILOOioiiO00OIl0lilllO ;
 wire [ 63: 0] Oo00IIIIoOIO0IL00llOoOioiollIOi00 ;
 wire [ 63: 0] OolIl0OOoiOlLioiloO0OolLOiIOolLLI ;
 wire [ 63: 0] OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ;
 wire [ 63: 0] O0lIi00lIl0iOlLilOloOIllllLLolooo ;
 wire [ 63: 0] OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ;
 wire [ 63: 0] O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ;
 wire [ 63: 0] OIoll0OLiliiLlIililii0oiII0Ol00lO ;
 wire [ 63: 0] Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ;
 wire [ 63: 0] OoOll0iOi0l0LiioLllOoliOoO00Lloil ;
 wire [ 63: 0] OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ;
 wire [ 63: 0] O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ;
 wire [ 63: 0] O0Il00oIILloI0IL0LiOO0i0lIiIoolio ;
 wire [ 63: 0] OI00OLIIi0LioLLLLllooOiOl0iolOO0I ;
 wire [ 63: 0] OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ;
 wire [ 63: 0] OOILLooOOlllIILoIiIioLIOI0LOiLiLI ;
 wire [ 63: 0] O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ;
 wire [ 63: 0] OOIoOIilLi0looLILloOOollIIIo0llLo ;
 wire [ 63: 0] O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ;
 wire [ 63: 0] OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ;
 wire [ 63: 0] OIIli0ilooIlOLI0lLO0Oi0IilILOolii ;
 wire [ 63: 0] OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ;
 wire [ 63: 0] OloILiOiLoIOOl0IoloOlI00Oollol0lL ;
 wire [ 63: 0] O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ;
 wire [ 63: 0] OI0ILilL0olIiOoL0lOiiooolOOllIIIL ;
 wire [ 63: 0] OIiIIlooOiolooLoI0iLi0loLiloiLOll ;
 wire [ 63: 0] OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ;
 wire [ 63: 0] OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ;
 wire [ 63: 0] OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ;
 wire [ 63: 0] OoOLolo0o0IOilOOLI0OoioLilIliI0lO ;
 wire [ 63: 0] OlOL0OLLooilLiOliIOIOOlIio00Oiili ;
 wire [ 63: 0] OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ;
 wire [ 63: 0] OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ;
 wire [ 63: 0] OlIliOioiio0LLoLl00i0liioIOI00iIi ;
 wire [ 63: 0] OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ;
 wire [ 63: 0] O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ;
 wire [ 63: 0] OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ;
 wire [ 63: 0] OLILoOooIiil0oIIolILIlLIioL0i0Iio ;
 wire [ 63: 0] O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ;
 wire [ 63: 0] Ol0LliIIIIiOOILo0ooioLolOOOololIo ;
 wire [ 63: 0] OIILiOiLOO0IILI0llIOoooi0oLiiOioO ;
 wire [ 63: 0] OiIoioILioOLl0io00oiOiO0liliOlOoO ;
 wire [ 63: 0] O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ;
 wire [ 63: 0] Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ;
 wire [ 63: 0] OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ;
 wire [ 63: 0] OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ;
 wire [ 63: 0] OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ;
 wire [ 63: 0] O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ;
 wire [ 31: 0] OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ;
 wire [ 31: 0] OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ;
 wire [ 31: 0] OIiLIoliOIilIl0O00Li00oIO0OlIiooo ;
 wire [ 31: 0] OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ;
 wire [ 31: 0] OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ;
 wire [ 31: 0] OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ;
 wire [ 31: 0] OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ;
 wire [ 31: 0] OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ;
 wire [ 31: 0] O0000LloLiliiLOoIi0iLiLli0iloOOLI ;
 wire [ 31: 0] OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ;
 wire [ 31: 0] OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ;
 wire [ 31: 0] OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ;
 wire [ 31: 0] Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ;
 wire [ 31: 0] O0o0OiliollLIi0IiLilIiOlLOOOLO00i ;
 wire [ 31: 0] OO0oolOlI0iloil0ooIolIioiol00I00I ;
 wire [ 31: 0] OLIoIliI0LI0liL0i0IIIiLloL000l0lO ;
 wire [ 31: 0] OO0iLILOLioOioLOoLIOlOlo0oOIollll ;
 wire [ 31: 0] OLOlLlooLIlL0IIiOilIiIooLloIioLOi ;
 wire [ 31: 0] OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ;
 wire [ 31: 0] OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ;
 wire [ 31: 0] O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ;
 wire [ 31: 0] OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ;
 wire [ 31: 0] OOI0llLoO0IOO000OilllLLLI0i0Iilil ;
 wire [ 31: 0] OlollLLLoL0iiI0lool0OOOOIiOoolioL ;
 wire [ 31: 0] OLOILIii00lILOLoLIIlOiioll0ilOLii ;
 wire [ 31: 0] OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ;
 wire [ 31: 0] O0OllOiIO00LliIOoLolo0loIiL0LiIlI ;
 wire [ 31: 0] Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ;
 wire [ 31: 0] OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ;
 wire [ 31: 0] OLIIl0o0liIOIooiOII0liO0oLllOI0oO ;
 wire [ 31: 0] Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ;
 wire [ 31: 0] OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ;
 wire [ 63: 0] OLli0lIO0lOO0OooILllIi00Lol00oili ;
 wire [ 63: 0] OOllI0oo0L0io0l0IoloioOii0oIioOi0 ;
 wire [ 63: 0] OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ;
 wire [ 63: 0] OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ;
 wire [ 63: 0] OoOOLol000OllOLI0LO0LO0LoIliO0iiL ;
 wire [ 63: 0] OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ;
 wire [ 63: 0] OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ;
 wire [ 63: 0] OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ;
 wire [ 63: 0] OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ;
 wire [ 63: 0] OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ;
 wire [ 63: 0] Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ;
 wire [ 63: 0] OiOoiILoiIiIIoll0loilLl00Ll00O0iL ;
 wire [ 63: 0] Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ;
 wire [ 63: 0] OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ;
 wire [ 63: 0] O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ;
 wire [ 63: 0] Oo00OloiOIoLi00Oo0ooiololoOoooLLO ;
 wire [ 63: 0] OI00OlLIOIiOOiIliIooII00LLLllLLOO ;
 wire [ 63: 0] OOlOiiLoIooll0L00oIIIoOIililiillo ;
 wire [ 63: 0] OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ;
 wire [ 63: 0] Oll00iO0Ol0IOLloLLilo0OliIloIiLli ;
 wire [ 63: 0] OIl0iolIOLOlLOloIoLoIo0OooLi000lO ;
 wire [ 63: 0] OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ;
 wire [ 63: 0] OOIOl00lliliioILLoiioolL0OLLoLo0i ;
 wire [ 63: 0] O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ;
 wire [ 63: 0] O0IlliiI0l00iOLL0oLilIILo00lLIolo ;
 wire [ 63: 0] OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ;
 wire [ 63: 0] OOOOLL0II0ioIiIIoLOolIOLIoLooIill ;
 wire [ 63: 0] OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ;
 wire [ 63: 0] OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ;
 wire [ 63: 0] OlOiOoL0i0i0L00OL00l00OOoL0OLILol ;
 wire [ 63: 0] OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ;
 wire [ 63: 0] Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ;
 wire [ 31: 0] Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ;
 wire [ 31: 0] OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ;
 wire [ 31: 0] O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ;
 wire [ 31: 0] OLLli0LLl0LlILOoi000iLoiiOOOLooLI ;
 wire [ 31: 0] OoIooi0LILolioIilliiol0I0iLoioIoi ;
 wire [ 31: 0] OILolilliOIlLILOoioLii0iI0lII0oil ;
 wire [ 31: 0] OOIilioOiLLoOIL0iLoILiLLliiio0LOl ;
 wire [ 31: 0] OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ;
 wire [ 31: 0] OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ;
 wire [ 31: 0] OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ;
 wire [ 31: 0] OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ;
 wire [ 31: 0] OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ;
 wire [ 31: 0] OioIoIoo0iIIlOilLlIoILioo0I0lo00o ;
 wire [ 31: 0] OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ;
 wire [ 31: 0] OLI00Il0O0lI0OoLI0oIloiOIiiILIill ;
 wire [ 31: 0] Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ;
 wire [ 31: 0] OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ;
 wire [ 31: 0] O0i000LoOoll00lolOOOOIO0Oio0LIO0o ;
 wire [ 31: 0] Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ;
 wire [ 31: 0] OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ;
 wire [ 31: 0] Oiio0oo000ioIO0llioIoLILlIlIOOloL ;
 wire [ 31: 0] OIooL0lILLIloiOOLiI0ilOIli0LOL000 ;
 wire [ 31: 0] OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ;
 wire [ 31: 0] OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ;
 wire [ 31: 0] OII0Iill0IOLO000li0iL0iLoiIoOoliL ;
 wire [ 31: 0] OOI0I0II0oOOO0LiLoO0I00LloOllilIl ;
 wire [ 31: 0] OOIioIlLoOL00lOliIIllL00illo0L00o ;
 wire [ 31: 0] OLiloooloollOoil0LlolLolOILlO00Ol ;
 wire [ 31: 0] OOilLILioilLIliOlOoilOOIolLLiLl0I ;
 wire [ 31: 0] OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ;
 wire [ 31: 0] OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ;
 wire [ 31: 0] OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ;
 wire OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ;
 wire Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ;
 wire Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ;
 wire OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ;
 wire OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ;
 wire OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ;
 wire O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ;
 wire OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ;
 wire OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ;
 wire OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ;
 wire OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ;
 wire OIlLiI0I0l0olLllLI0LliOOlllliLL0i ;
 wire O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ;
 wire OOIILlIiIOiOIi0o0li0lolol0LIoOliI ;
 wire OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ;
 wire Ollil0L0OlO0loio0OLiLILo0OioO0iOO ;
 wire O0L0O0ioooOOiLLlLLOLiioooILolII0o ;
 wire OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ;
 wire OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ;
 wire OLllIIIO0oIlllOo00LILooILo0io0o00 ;
 wire OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ;
 wire O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ;
 wire OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ;
 wire OllloLIILloiiiOill0lOLooilli0Llii ;
 wire OoIL0ll0llIOoI0IoIioiILILllLLOOOL ;
 wire OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ;
 wire OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ;
 wire O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ;
 wire OiOo0O0ooiioi00lloILL0oLLoILOiLiO ;
 wire OlLILiOolLl0ioiLiLlILiILLlIOllloI ;
 wire OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ;
 wire O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ;
 wire [ 15: 0] OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ;
 wire OOooLlloIiioOOO0LLILl0liiillLILol ;
 wire [31:0] OoOi0O0oOoL0looLo0IoOllOOILiLooLl ;
 wire [31:0] OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO ;
 wire [31:0] OLlOiiLlLoolliOiO0i0lOloio0L0oL00 ;
 wire [31:0] OilOI0i0lloo0Lll000I0OIoIOI0lioiO ;
 wire [31:0] OlooiiLooL0L00oIIiioLloiIolOoOlLo ;
 wire [31:0] OLo0LOlILllLILOIiiiL0LIlLIoLlO0II ;
 wire [31:0] OiiOioOIO00LOOLilooiooo0olO0illo0 ;
 wire [31:0] OLl0LoLoii00oiOOoilollii000iIOlOI ;
 wire [31:0] OLlil0000Oiil0IOOLiloIlliOoLLol0L ;
 wire [31:0] OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI ;
 wire [31:0] OO0OOILiO000LOILL0OllLi0l0oliLOo0 ;
 wire [31:0] OLiLllIIIlo0llILiLloLOoooOLOilI0l ;
 wire [31:0] Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl ;
 wire [31:0] OiL0IiiliiioOOLliLiiLILlIOloOLL0L ;
 wire [31:0] OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi ;
 wire [31:0] OllLOLiIilI0oili000OiLilLioIOoIl0 ;
 wire [31:0] OOooI0loOL0iiOIoOili0OOOLLiiIiLOl ;
 wire [31:0] OLIIiIIIOILl0loi0lO0IiOoolLIloi00 ;
 wire [31:0] OoOillIILLoLoOioLloli0OLILlIOOoLo ;
 wire [31:0] OlOlO00LLloOiOolOiOLOIiloLil0L0LI ;
 wire [31:0] OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO ;
 wire [31:0] OlOLIILoL0ll0oooOo0OIoLoOoiLIolol ;
 wire [31:0] OIlLOILiLLo0ol0OLlI0IILilILLLlILO ;
 wire [31:0] O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i ;
 wire [31:0] Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL ;
 wire [31:0] OOiIlillllLOI0oOOoILlol0ILoIoOLil ;
 wire [31:0] OOIiO0olO0OLlo0liIoiOioiIO00oOIiL ;
 wire [31:0] O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 ;
 wire [31:0] OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l ;
 wire [31:0] OlolLlliLo0O0l0lOOolL0ioI0O0Li00l ;
 wire [31:0] Oo0oI0oLOLlloloiiLIIol0LilOlOIliI ;
 wire [31:0] OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo ;
 wire [31:0] OoiLlL0oiiIloLOoloIL0oLii00IIIoII ;
 wire [31:0] Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ;
 wire [15:0] Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 wire [31:0] OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ;
 wire [31:0] OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ;
 wire O0OlOIIOOIOIioo00liool0iIiI0I0Lll ;
 wire [ 3:0] O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii ;
 wire OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l ;
 wire OIiOIl0O0OLllloOl0oOoLoIllIL0illO ;
 wire [63:0] Oi0loi0OllIlIoI0ILloIllILIO0IIo0I ;
 wire [ 2:0] OoLOIol0OLIIiloO0oLoiliOl0LilIolI ;
 wire [15:0] OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i ;
 wire [15:0] OOloOOOOiILOioIlIOO0oILilOLLL00OO;
 wire [31:0] OOIlIOO0IL0OoLli0IoliIioOOlIILlii ;
 wire OoI0IoiILOOLILioiioIOoOLioiiOlIio ;
 wire OioOlll0OooLLL0IIIIIli0ollooo0L0L ;
 wire [15:0] OooOLOOliIlIOlio00OO0oloLoOi0lliO ;
 wire [15:0] OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI ;
 wire [15:0] OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL ;
 wire [15:0] Oo0OiL0Lll000LlioLiooLOLloiLiliii ;
 wire [15:0] OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI ;
 wire [15:0] OioiIooIlil0liIiOIi0lLLIllOioioli ;
 wire [15:0] OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 ;
 wire [15:0] OlLloLOlOi0iIiLIlOlLio000LLOLILli ;
 wire [15:0] OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 ;
 wire [15:0] OOlILOLoilIOloioiIoOLI0L0ooLO0Lll ;
 wire [15:0] OolOlIOiIIoII0ll0IllLoOiIllIilOoO ;
 wire [15:0] OOIiiol0IOILiLloOLiLOIIlIIolooOIO ;
 wire [15:0] OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO ;
 wire [15:0] OILili00ILILlO0LIoLlll0oliLio0liL ;
 wire [15:0] OoILoooiioLLiIIIoiIoiOIO0OllIlIlL ;
 wire [15:0] OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO ;
 wire [15:0] OIiiiIlLolLIoIioOoOolloi0L0loLoIL ;
 wire [15:0] OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO ;
 wire [15:0] O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II ;
 wire [15:0] OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO ;
 wire [15:0] OOlO0o0i0Io0IOllLoIloiioiliOOlIII ;
 wire [15:0] OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I ;
 wire [15:0] O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 ;
 wire [15:0] OlOlLO00i0Oiooo0lLollo0IILIlLO0OI ;
 wire [15:0] OLLliI0IiOiollllIOOLL0oL0IlllO0oI ;
 wire [15:0] OLO00iLliol0LLIOOIIO0IiLIllO0IL0O ;
 wire [15:0] O0OII0Ili0ilol00OLOLoiOl0OlLo0liO ;
 wire [15:0] OOL0lolilI0oIloIoIIILooo0lOLOlolI ;
 wire [15:0] OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll ;
 wire [15:0] OIO00IOolLoOoOL0ILI00i0olI0IiiOOo ;
 wire [15:0] OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO ;
 wire [15:0] OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 ;
 wire [15:0] OIoiIlOo00oL0iL0o0iooollLlilLoIIo ;
 wire O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ;
 output [3:0] OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI ;
 output OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 ;
 output [5:0] OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI ;
 output OilOOo00lLiOOoiO0ii0oo0oOliOollii ;
 output [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 output [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 wire [3:0] OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI ;
 wire OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 ;
 wire [5:0] OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI ;
 wire OilOOo00lLiOOoiO0ii0oo0oOliOollii ;
 wire [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 wire [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 wire [15:0] O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ;
 wire OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 wire [ 15:0] OILIloOoilLIL00IIOoOilLOO0L0iiIOO ;
 wire [ 31:0] O0oLLi0Ill00l0lioiLioiooIllloIiIl ;
 wire OOiiOOiio0liOLLo00IOILoIi0lIli0I0 ;
 wire Oo0LOIoiLLilIiOlLiIlLOi0OOLOooO0i ;
 wire O0iIiiLOl0llolLOO0iliI0L00LoliL0O ;
 wire O0IOlOo0oLillLIiLli0LiI0oIIlo0Loo ;
 wire OiLiiLIlIO0O0oIliIlLiOlolOlIll0LO ;
 wire OLoIIlo0lILOLILillIOOilOIilLillO0 ;
 wire OIiiOiO0i00Li0OOl0oo0IOLILioo0L0l ;
 wire OIIOOLloiL0IoIlLliLolILlIiOIILiOI ;
 wire OLl0L0IIoOoIi0iiIO000IIIiLoi0IiLo ;
 wire O00LLILiIoI00LOOoiLlI0oLIiiL0OOI0 ;
 wire Olo0ILLoliIOlOOo0OIo0Lllo0oiLOIlI ;
 wire OLioiooIL0o0oiILiolOLi0Ll0iOoiOII ;
 wire O0lIO0LlOooLILO0iLlLLIiIlLiiolOiO ;
 wire OllooIiliLOIOoIoLoOII0LLLii0O0IIL ;
 wire OlILIiOOIOlLiLiLiiLO0LI0I0LliL0oL ;
 wire OLIIiiLOlO0LLLiOlO0O0Oo0LOLLiILoI ;
 wire OiOooooIliLiLL00i0loL00ol0LooI0II ;
 wire Oi0ilOLi0LOOoO00Oi0LiIOo0I0oLilIO ;
 wire OlIOlOillOlO0ol0iolIlLOiooOio0LOi ;
 wire OIl0oIiIIiLiIiLOiOOLOI0lOOOIIiIoo ;
 wire O0oLiLiLlOlIIiLoLiLIiLL0l0oI0iIlO ;
 wire O0IL0iiIilolIlIiLIIIIOOiLOoOoloLL ;
 wire O0ILooiI0L00OoOoLlL0i0OooLOolooiO ;
 wire OO0ooiOliiL0l0OoiiloO0oLIIIioII0L ;
 wire O0iilOLolIOOlILi0iI0LLlLloiLO0L0O ;
 wire OIILI00Loo0ooOiOL000Ilo00ool0I0oo ;
 wire OOooo0i0LloOLo00OIOIllLLiILOLLll0 ;
 wire OlLlL0ilOI0II0l0ILLIlIOLOoI0LiLIi ;
 wire O0Ll0LoIi00OO0iolo0ILiolI0LOolooi ;
 wire Ool0o0OoOlOiL00i00O0iloIO0Lo00oOI ;
 wire OIlOi0LL0LOLOLLL0LIIio0LLliiIoilo ;
 wire OilOOiiLIo0ooi0OLoliio0iooIooil0o ;
 wire [31:0] Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 0] = OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 1] = Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 2] = Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 3] = OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 4] = OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 5] = OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 6] = O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 7] = OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 8] = OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 9] = OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[10] = OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[11] = OIlLiI0I0l0olLllLI0LliOOlllliLL0i ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[12] = O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[13] = OOIILlIiIOiOIi0o0li0lolol0LIoOliI ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[14] = OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15] = Ollil0L0OlO0loio0OLiLILo0OioO0iOO ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[16] = O0L0O0ioooOOiLLlLLOLiioooILolII0o ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[17] = OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[18] = OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[19] = OLllIIIO0oIlllOo00LILooILo0io0o00 ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[20] = OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[21] = O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[22] = OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23] = OllloLIILloiiiOill0lOLooilli0Llii ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[24] = OoIL0ll0llIOoI0IoIioiILILllLLOOOL ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[25] = OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[26] = OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[27] = O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[28] = OiOo0O0ooiioi00lloILL0oLLoILOiLiO ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[29] = OlLILiOolLl0ioiLiLlILiILLlIOllloI ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[30] = OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31] = O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ;
 assign OOooLlloIiioOOO0LLILl0liiillLILol = OOiiOOiio0liOLLo00IOILoIi0lIli0I0 || Oo0LOIoiLLilIiOlLiIlLOi0OOLOooO0i || O0iIiiLOl0llolLOO0iliI0L00LoliL0O || O0IOlOo0oLillLIiLli0LiI0oIIlo0Loo || OiLiiLIlIO0O0oIliIlLiOlolOlIll0LO || OLoIIlo0lILOLILillIOOilOIilLillO0 || OIiiOiO0i00Li0OOl0oo0IOLILioo0L0l || OIIOOLloiL0IoIlLliLolILlIiOIILiOI || OLl0L0IIoOoIi0iiIO000IIIiLoi0IiLo || O00LLILiIoI00LOOoiLlI0oLIiiL0OOI0 || Olo0ILLoliIOlOOo0OIo0Lllo0oiLOIlI || OLioiooIL0o0oiILiolOLi0Ll0iOoiOII || O0lIO0LlOooLILO0iLlLLIiIlLiiolOiO || OllooIiliLOIOoIoLoOII0LLLii0O0IIL || OlILIiOOIOlLiLiLiiLO0LI0I0LliL0oL || OLIIiiLOlO0LLLiOlO0O0Oo0LOLLiILoI || OiOooooIliLiLL00i0loL00ol0LooI0II || Oi0ilOLi0LOOoO00Oi0LiIOo0I0oLilIO || OlIOlOillOlO0ol0iolIlLOiooOio0LOi || OIl0oIiIIiLiIiLOiOOLOI0lOOOIIiIoo || O0oLiLiLlOlIIiLoLiLIiLL0l0oI0iIlO || O0IL0iiIilolIlIiLIIIIOOiLOoOoloLL || O0ILooiI0L00OoOoLlL0i0OooLOolooiO || OO0ooiOliiL0l0OoiiloO0oLIIIioII0L || O0iilOLolIOOlILi0iI0LLlLloiLO0L0O || OIILI00Loo0ooOiOL000Ilo00ool0I0oo || OOooo0i0LloOLo00OIOIllLLiILOLLll0 || OlLlL0ilOI0II0l0ILLIlIOLOoI0LiLIi || O0Ll0LoIi00OO0iolo0ILiolI0LOolooi || Ool0o0OoOlOiL00i00O0iloIO0Lo00oOI || OIlOi0LL0LOLOLLL0LIIio0LLliiIoilo || OilOOiiLIo0ooi0OLoliio0iooIooil0o ;
 OiI00lI0lL0IoLLLlLoioLlOIOOiOiiIi OiI00lI0lL0IoLLLlLoioLlOIOOiOiiIi ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L (Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L), .OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl (OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl), .OoIolioOL0iLLOLloI00iIILLiiL0Ooil(OoIolioOL0iLLOLloI00iIILLiiL0Ooil), .Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 ) , .OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI (OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI), .OLOILlOloOoi0OO0oLOOlo0iiIoioilL0(OLOILlOloOoi0OO0oLOOlo0iiIoioilL0), .OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI(OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI) , .OilOOo00lLiOOoiO0ii0oo0oOliOollii (OilOOo00lLiOOoiO0ii0oo0oOliOollii) , .OOLIiil0IlIllLollIl0LIilliOI0iolo (OOLIiil0IlIllLollIl0LIilliOI0iolo ), .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl ), .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ), .O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo (O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ), .OILIloOoilLIL00IIOoOilLOO0L0iiIOO (OILIloOoilLIL00IIOoOilLOO0L0iiIOO), .O0oLLi0Ill00l0lioiLioiooIllloIiIl (O0oLLi0Ill00l0lioiLioiooIllloIiIl), .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 (OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ), .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ), .OLo0oiiL0ooIliO0I0illLoILiiIoIoOI (OLo0oiiL0ooIliO0I0illLoILiiIoIoOI), .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi), .OoiloolOiOIoIOolLiOl0OlOiOli0oOOl (OoiloolOiOIoIOolLiOl0OlOiOli0oOOl), .OillLliLoolOIiiiILoOILOIloo000iLI (OillLliLoolOIiiiILoOILOIloo000iLI), .OlLOLoI0iIOLloliOllILlOoIiioOli0L (OlLOLoI0iIOLloliOllILlOoIiioOli0L), .Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ), .O0Loo0iiI0OlLOlOIiILOooOOlIoioOli (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ), .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl), .OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO (OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO), .OLlOiiLlLoolliOiO0i0lOloio0L0oL00 (OLlOiiLlLoolliOiO0i0lOloio0L0oL00), .OilOI0i0lloo0Lll000I0OIoIOI0lioiO (OilOI0i0lloo0Lll000I0OIoIOI0lioiO), .OlooiiLooL0L00oIIiioLloiIolOoOlLo (OlooiiLooL0L00oIIiioLloiIolOoOlLo), .OLo0LOlILllLILOIiiiL0LIlLIoLlO0II (OLo0LOlILllLILOIiiiL0LIlLIoLlO0II), .OiiOioOIO00LOOLilooiooo0olO0illo0 (OiiOioOIO00LOOLilooiooo0olO0illo0), .OLl0LoLoii00oiOOoilollii000iIOlOI (OLl0LoLoii00oiOOoilollii000iIOlOI), .OLlil0000Oiil0IOOLiloIlliOoLLol0L (OLlil0000Oiil0IOOLiloIlliOoLLol0L), .OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI (OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI), .OO0OOILiO000LOILL0OllLi0l0oliLOo0 (OO0OOILiO000LOILL0OllLi0l0oliLOo0), .OLiLllIIIlo0llILiLloLOoooOLOilI0l (OLiLllIIIlo0llILiLloLOoooOLOilI0l), .Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl (Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl), .OiL0IiiliiioOOLliLiiLILlIOloOLL0L (OiL0IiiliiioOOLliLiiLILlIOloOLL0L), .OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi (OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi), .OllLOLiIilI0oili000OiLilLioIOoIl0 (OllLOLiIilI0oili000OiLilLioIOoIl0), .OOooI0loOL0iiOIoOili0OOOLLiiIiLOl (OOooI0loOL0iiOIoOili0OOOLLiiIiLOl), .OLIIiIIIOILl0loi0lO0IiOoolLIloi00 (OLIIiIIIOILl0loi0lO0IiOoolLIloi00), .OoOillIILLoLoOioLloli0OLILlIOOoLo (OoOillIILLoLoOioLloli0OLILlIOOoLo), .OlOlO00LLloOiOolOiOLOIiloLil0L0LI (OlOlO00LLloOiOolOiOLOIiloLil0L0LI), .OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO (OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO), .OlOLIILoL0ll0oooOo0OIoLoOoiLIolol (OlOLIILoL0ll0oooOo0OIoLoOoiLIolol), .OIlLOILiLLo0ol0OLlI0IILilILLLlILO (OIlLOILiLLo0ol0OLlI0IILilILLLlILO), .O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i (O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i), .Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL (Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL), .OOiIlillllLOI0oOOoILlol0ILoIoOLil (OOiIlillllLOI0oOOoILlol0ILoIoOLil), .OOIiO0olO0OLlo0liIoiOioiIO00oOIiL (OOIiO0olO0OLlo0liIoiOioiIO00oOIiL), .O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 (O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0), .OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l (OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l), .OlolLlliLo0O0l0lOOolL0ioI0O0Li00l (OlolLlliLo0O0l0lOOolL0ioI0O0Li00l), .Oo0oI0oLOLlloloiiLIIol0LilOlOIliI (Oo0oI0oLOLlloloiiLIIol0LilOlOIliI), .OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo (OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo), .OoiLlL0oiiIloLOoloIL0oLii00IIIoII (OoiLlL0oiiIloLOoloIL0oLii00IIIoII), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO (Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ), .OOllOo00o0IlooI0l0io0O00l0OIoiILO (OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ), .OOiiILlloiOoI0OlilIOoiiLOOLol0IoI (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ), .OiiLOILl0iLi0L0ilIIoooLLIoliIIIlO ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OOOLiLOilooIi0Iio00ilILoLIILOoOoI ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( O0OlOIIOOIOIioo00liool0iIiI0I0Lll ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OIiOIl0O0OLllloOl0oOoLoIllIL0illO ) , .OL0O0IIio0loL0L0Il0li0i00lliIoOOI ( OL0O0IIio0loL0L0Il0li0i00lliIoOOI ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( Oi0loi0OllIlIoI0ILloIllILIO0IIo0I ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OoLOIol0OLIIiloO0oLoiliOl0LilIolI ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i ) , .OilOOioILlOIIOL0iioIOIi0oloooOoLl ( OOloOOOOiILOioIlIOO0oILilOLLL00OO ) , .OI00OiLolooiIIiiILoIliO0O0loolIlI ( OioOlll0OooLLL0IIIIIli0ollooo0L0L ) , .OOL0o0i0Llo0IiiLlO00oliOILLI00Ool ( OOIlIOO0IL0OoLli0IoliIioOOlIILlii ) , .OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ( OooOLOOliIlIOlio00OO0oloLoOi0lliO ) , .OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo (OoI0IoiILOOLILioiioIOoOLioiiOlIio ) , .OIloLiiOL00oilLo0iiILoOOll0lIlIlO ( OIloLiiOL00oilLo0iiILoOOll0lIlIlO ) , .Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ( Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ) , .O0oill0llILOilo0i0LIoOLIoolL0Il0o (O0oill0llILOilo0i0LIoOLIoolL0Il0o ) , .OlliILlLOilOl0LO0O0OilooiIIiOi0Ll (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) , .OOLoL0looIOoioIoOooIoLIiIiLiLoiOl (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) , .OIoIooIolOilIOlooOlOIIOoilLioOIIO (OIoIooIolOilIOlooOlOIIOoilLioOIIO ) , .OiL0LolLLIOlliloII00llOil0oIlOiIo (OiL0LolLLIOlliloII00llOil0oIlOiIo ) , .O0llIOIliLOO0iiOoO0OO0lIOloLoII0I (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ) , .OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL ) , .OilOIloOO0LiLoIL0IIILoIi0Loilll0I ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I ) , .Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ) , .OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ) , .OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ( OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ) , .OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ( OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ) , .OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ( OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ) , .OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ( OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ) , .OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ( OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ) , .OiooiLLioLLL0lII00ol0oIOllLlOiLlL ( OiooiLLioLLL0lII00ol0oIOllLlOiLlL ) , .OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ( OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ) , .O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ( O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ) , .Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ( Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ) , .O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ( O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ) , .OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ( OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ) , .OilLIO0lI0LO0LolOOilILl0oiIlolOlo ( OilLIO0lI0LO0LolOOilILl0oiIlolOlo ) , .OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ( OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ) , .OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ( OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ) , .OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ( OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ) , .OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ( OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ) , .OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ( OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ) , .OIoliiOo0i000ooilOOLOiil0LlLiOoLo ( OIoliiOo0i000ooilOOLOiil0LlLiOoLo ) , .Oo00OlooOo0io0OoIloiioLiOlL0llio0 ( Oo00OlooOo0io0OoIloiioLiOlL0llio0 ) , .OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ( OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ) , .OOoOoILioOoIlIoLliOLOOi0io0IlLolo ( OOoOoILioOoIlIoLliOLOOi0io0IlLolo ) , .OiLllooo0Li0lioiolLi0ILIoLOliil0I ( OiLllooo0Li0lioiolLi0ILIoLOliil0I ) , .OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ( OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ) , .OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ( OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ) , .OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ( OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ) , .OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ( OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ) , .OLL0OiLILloil0IoOlLIIloLIiIlllLil ( OLL0OiLILloil0IoOlLIIloLIiIlllLil ) , .OILI0LLillilOlllLil0ioLoIiliOoLLo ( OILI0LLillilOlllLil0ioLoIiliOoLLo ) , .OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ( OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ) , .OoIloII0oLiOLOLIllOL0iOoooOliOIii ( OoIloII0oLiOLOLIllOL0iOoooOliOIii ) , .Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ( Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ) , .OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ( OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ) , .OO0liOO0iOOIioool0OoLliiiI0l0ilOo ( OO0liOO0iOOIioool0OoLliiiI0l0ilOo ) , .OiIOLi00lOILlOOL0oLLloL0io0LoIoOL (OiIOLi00lOILlOOL0oLLloL0io0LoIoOL) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OOooLlloIiioOOO0LLILl0liiillLILol ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OloliIooiiLI0IIlOiL0LLlioILLllL0L ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OioILlIiO0000OoolooO00loIOIloLIoI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLOl0000OLooLIIo0lIOIOI0lILioolOl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OoIolLlOIIoIoi00lloLlIoI0lo0iILol ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOIIloOlOILliIOILOIOiIlooIOOIL0oO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( O0liLooiLliIoLOllliIlo0ILo0I0oOOl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0i00oOl00OoIIOIil0LLOi0looIOIL00 ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OoOil0iLoliioLioOOilL0OlOO0IIOoI0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[0] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[0] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[0] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[0] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[0] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[0] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[0] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OOiiOOiio0liOLLo00IOILoIi0lIli0I0 ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OoolLolOioLILoOIII00LIOli00LIlloi ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OOOooLlOLO0iOOOLi00oIiloILlooOLIO ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OioLioLloIiilLLoOlIoiLIO0IOoiLoll ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OIiO0OLioLiIOIIiLoiLooI00I0olI00O ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OOOo0I0LlloiIl0i0il0OLiOlooOOolil ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OLlOlii00IoIl00oIioIiIool0lLiOoLo ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OIollo0oLlLiI0IILOO00illIILLIoo0o ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OLli0lIO0lOO0OooILllIi00Lol00oili ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OO0OIilooOLiLlollOiOLLo0LOOll0oo0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLlOiiLlLoolliOiO0i0lOloio0L0oL00 ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[1] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[1] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[1] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[1] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[1] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[1] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[1] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( Oo0LOIoiLLilIiOlLiIlLOi0OOLOooO0i ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OOIolooo0Oi00io00lIiiOiiLIliliOio ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OoI00LooIIlIIlIOOLIoloilI0OoIILLi ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OOIoOIilLi0looLILloOOollIIIo0llLo ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOllI0oo0L0io0l0IoloioOii0oIioOi0 ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII Olili0IOOooLOiOO0I00Oolil0oloOLl0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OilOI0i0lloo0Lll000I0OIoIOI0lioiO ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[2] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[2] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[2] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[2] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[2] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[2] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[2] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0iIiiLOl0llolLOO0iliI0L00LoliL0O ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( Oo0OiL0Lll000LlioLiooLOLloiLiliii ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( O0oLiillllLOiLilOoI000iOLoiL0L0LO ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OI0ioOlloiIio0oiOloi0lioiILoollLl ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OlIloooO00OIL0L0iIili0iOOoiLI0oiI ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OolIilIL0iooOLllOLloloOIlLIiOoLo0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O0lIOiilLOiIOollILlioiiOOiiLOO00i ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OIiLIoliOIilIl0O00Li00oIO0OlIiooo ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOiiiLlilOoOoOOOOoL0ii0LOLOiO0l00 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OlooiiLooL0L00oIIiioLloiIolOoOlLo ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[3] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[3] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[3] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[3] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[3] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[3] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[3] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0IOlOo0oLillLIiLli0LiI0oIIlo0Loo ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OOoL0lOOloLLOLOILLLOolliIll0oOOoO ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( Ol000OloII0LlIII00IIOIlOiioOo0Iii ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OLLli0LLl0LlILOoi000iLoiiOOOLooLI ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OilILLloOiOliioI00oOLililLO0oL0iO ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLo0LOlILllLILOIiiiL0LIlLIoLlO0II ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[4] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[4] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[4] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[4] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[4] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[4] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[4] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OiLiiLIlIO0O0oIliIlLiOlolOlIll0LO ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OioiIooIlil0liIiOIi0lLLIllOioioli ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OoooIiooOl0i0oliO0lio0IOo0iIILLLi ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OoOlILlliliiOI0OLLoOOl0000iIo0IIo ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLolLol0lLIIlIillI000oIlilLLloOii ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OO0O0oOlliIoIOlooIO0lOLolIilLllIO ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( O00I0iOoILll0oILl0ILloii0LIIOOiIO ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OlolloloolOo0o0LLLIl00Li0iiLl00ol ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OIIli0ilooIlOLI0lLO0Oi0IilILOolii ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OoOOLol000OllOLI0LO0LO0LoIliO0iiL ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OoIooi0LILolioIilliiol0I0iLoioIoi ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOOI0oOoioii0Lli0o0lL0OLoiLiOII0i ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OiiOioOIO00LOOLilooiooo0olO0illo0 ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[5] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[5] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[5] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[5] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[5] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[5] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[5] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OiooiLLioLLL0lII00ol0oIOllLlOiLlL ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OLoIIlo0lILOLILillIOOilOIilLillO0 ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLlLoL0lO0oOIOolIIoiILIO0oOilooll ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O0iI0Lil0liLOLiILLOoilII0LII0iolO ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OLLloO00IliLiLLlLloLloO0liOoIIOOI ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OO00IIiOlOioiOLIiIloilLII0lLL0OOi ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOLIlLlLIloIOoooilolooLloIi0OiiIi ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OILolilliOIlLILOoioLii0iI0lII0oil ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOoLlIiOo0lLilILLiiOOOIillLiO0ol0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLl0LoLoii00oiOOoilollii000iIOlOI ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[6] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[6] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[6] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[6] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[6] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[6] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[6] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OIiiOiO0i00Li0OOl0oo0IOLILioo0L0l ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OlLloLOlOi0iIiLIlOlLio000LLOLILli ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OoLLliL00LLoooll00ooiLolOliOO0lLI ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O00loOoIIlII0OOo0lio00iOOOolLiIiO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OiiOIoolI0LioIo0IlL0lOllILIOOiIio ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OoIooolIllLIIolLII0IiLLiiOlOOIIOO ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OLL0i00LllLlio0oLOLooIL0ilLLllil0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OOiOiOIIoOii0oOLlI0OliIi0liioLLII ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OlOl0iOIioolOiill0OLOloOoLiIlllol ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OloILiOiLoIOOl0IoloOlI00Oollol0lL ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OOIilioOiLLoOIL0iLoILiLLliiio0LOl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OiiI0iLOloILO0LlOLLOOOOl0L0l0l0Oo ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLlil0000Oiil0IOOLiloIlliOoLLol0L ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[7] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[7] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[7] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[7] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[7] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[7] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[7] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OIIOOLloiL0IoIlLliLolILlIiOIILiOI ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( O0li0llLIi0oIo0IilLLooLILolLIOOoo ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OioIOIo0IllIo0OILLlli0LOOl00lioII ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OLOoO0oILOiOlioILlooiILlll0iiiL0O ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[8] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[8] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[8] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[8] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[8] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[8] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[8] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OLl0L0IIoOoIi0iiIO000IIIiLoi0IiLo ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OOlILOLoilIOloioiIoOLI0L0ooLO0Lll ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0il0OIIioo0IoL0OI0llOiLiLioill0i ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( O0lioOi00lO0IL00IoLLILolIlli00LiI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OioOlIooLl0IL0LiioIlILIolO0o0ii0l ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OI0ILilL0olIiOoL0lOiiooolOOllIIIL ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( O0000LloLiliiLOoIi0iLiLli0iloOOLI ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII O0liio0IOOlOIo0IoiiLLooLO0lLiL0Oo ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OO0OOILiO000LOILL0OllLi0l0oliLOo0 ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[9] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[9] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[9] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[9] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[9] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[9] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[9] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O00LLILiIoI00LOOoiLlI0oLIiiL0OOI0 ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OolOlIOiIIoII0ll0IllLoOiIllIilOoO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OIO0IIi0OIooOiLOIII0lLolililiOIll ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OioilLoll0OiiOooiLiIOiL0LiilILII0 ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OLoli0Li0i0oO0olOOilIliIio0LOoIIO ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OLLOoOIo0oiL0IOOO0lill0iloILllIOO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OIILOOOOIOl00OoIollioiiliIilolLLl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OiooooLLoI0OLilIIil0ilooLo0OIloLl ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OiLiiLILIoLilioiLolliOl0LI00LLil0 ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( Oloo0IIooolliliLOLoLoL0oI0LOliLlL ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OIiIIlooOiolooLoI0iLi0loLiloiLOll ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OO0lO0o0L0oioloiiI0o0lILILLoLiLlo ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLiLllIIIlo0llILiLloLOoooOLOilI0l ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[10] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[10] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[10] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[10] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[10] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[10] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( Olo0ILLoliIOlOOo0OIo0Lllo0oiLOIlI ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OOIiiol0IOILiLloOLiLOIIlIIolooOIO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( Ol0OLoIiI0OloLIlillLOloLioIIL0III ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OiILooool0OiolIOIIlO0LiOliIiIL0Ii ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OlLiiOLII0io0OLOOiIiiO0IIililoolo ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLlolloLliiLO0IlIlLo0lIiiloL00OOL ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O00oIiiOLOoilolOol0OIIOII00lllOIo ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OLiIOloOILlLO0IlooI0lo0OI0OOIiooi ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[11] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[11] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[11] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[11] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[11] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[11] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OilLIO0lI0LO0LolOOilILl0oiIlolOlo ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OLioiooIL0o0oiILiolOLi0Ll0iOoiOII ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLi0ooOo0OlIllLOILllLL00lL00Liii0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OOOLilOolI0LILLIoloIiO00OiIiLiiIo ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OlLi0LOI0LoLioI0loilIlo00iliILIoi ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OiOoiILoiIiIIoll0loilLl00Ll00O0iL ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OIlLiI0I0l0olLllLI0LliOOlllliLL0i ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OilIoIiOlOIioOOi0oI0ILolooIioiILI ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OiL0IiiliiioOOLliLiiLILlIOloOLL0L ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[12] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[12] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[12] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[12] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[12] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[12] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0lIO0LlOooLILO0iLlLLIiIlLiiolOiO ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OILili00ILILlO0LIoLlll0oliLio0liL ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OO0OOoLL0O0OOOllioILi0liilLLloiLO ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OlLlliliOioioOIoiLOIOiOoiiioIOLOO ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OliliILl0LLiioool00L00LoLLILio0lO ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OLioIOLOILilililoO0ililOi0oiIoo0o ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OioIoIoo0iIIlOilLlIoILioo0I0lo00o ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OoLllLoOIIoolLlio0IIOIOo0i0LIIilL ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[13] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[13] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[13] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[13] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[13] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[13] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OllooIiliLOIOoIoLoOII0LLLii0O0IIL ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OoILoooiioLLiIIIoiIoiOIO0OllIlIlL ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OoLiLLooILIo0iol0OIoliLi0iiioiIlI ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OI0ool0i0ollOOoloL00L0LlLIO0LIliI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( Oo0loliLllliloIiliOi0lILloLI0ILlO ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( Ooi0OL0i0IioliooLiI00OoiL00looOIL ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OoOLolo0o0IOilOOLI0OoioLilIliI0lO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( O0o0OiliollLIi0IiLilIiOlLOOOLO00i ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OOIILlIiIOiOIi0o0li0lolol0LIoOliI ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII O0i0LiiiiLooLIi0IlOILiIIo00lO0IOL ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OllLOLiIilI0oili000OiLilLioIOoIl0 ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[14] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[14] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[14] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[14] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[14] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[14] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OlILIiOOIOlLiLiLiiLO0LI0I0LliL0oL ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OOIlIio0iILll00lliIIioiIiOLlLLi00 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OlIollIiLi0IlLiolloLOOL000Oo0l0II ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OiiooiLLOL0iiO0oILoOlLoololiIIo0o ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OL0Lio0lIililolilllOL0Li0lIi0I0LI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OolL0oo00LOo0LOoLiILllLo0loOoIiii ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OIOIOlilIolIlLOLlLlll0IiOIiILiOol ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OiloLLIlO00Il0oo0io0Iilliiil0OolO ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( O0oOL0illOloooo0ioIiOLOooLILllLl0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OlOL0OLLooilLiOliIOIOOlIio00Oiili ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OO0oolOlI0iloil0ooIolIioiol00I00I ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OLI00Il0O0lI0OoLI0oIloiOIiiILIill ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OiOIioILlIOlOi0IlIllOlOOlliIOIo0l ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OOooI0loOL0iiOIoOili0OOOLLiiIiLOl ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[15] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[15] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[15] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[15] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[15] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[15] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OLIIiiLOlO0LLLiOlO0O0Oo0LOLLiILoI ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OIiiiIlLolLIoIioOoOolloi0L0loLoIL ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOoLol0oioL0looOlO0io0oIillil0iI0 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( O0oilLoOiOiLLi0Li0lLOIooIiliILlii ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OLiILioillIololIOILoOLlI0LILLliIL ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OoOOillllIiloIOIILO0lL0LIl0iOlIII ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OLIoIliI0LI0liL0i0IIIiLloL000l0lO ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( Oo00OloiOIoLi00Oo0ooiololoOoooLLO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( Ollil0L0OlO0loio0OLiLILo0OioO0iOO ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OIoO0lIIOlol0LLilo0LOiLlIOiiOo0LL ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OLIIiIIIOILl0loi0lO0IiOoolLIloi00 ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[16] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[16] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[16] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[16] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[16] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[16] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OiOooooIliLiLL00i0loL00ol0LooI0II ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLio000LoL0lOol0oIiLlILLIlOLLOIlO ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OILIi00LOILOoLIiLloLiLIolliOoooIo ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OioilI0Oo0oOil0lIioiILIOLLLOLLioO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OI0L0iIOilOi0LlILL0l0liiiil0lOIii ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OlIIioIIlILoli0oIiIl0l0IlOlloooll ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OIOO0oiiIiiOILOOioiiO00OIl0lilllO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OO0iLILOLioOioLOoLIOlOlo0oOIollll ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OI00OlLIOIiOOiIliIooII00LLLllLLOO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0L0O0ioooOOiLLlLLOLiioooILolII0o ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII Oool0lLlloOIOlLOlo0iOIliIloo0i0IL ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OoOillIILLoLoOioLloli0OLILlIOOoLo ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[17] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[17] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[17] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[17] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[17] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[17] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OIoliiOo0i000ooilOOLOiil0LlLiOoLo ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( Oi0ilOLi0LOOoO00Oi0LiIOo0I0oLilIO ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OoiiooOo00OI0O0loiolLOLioIOiI0LoI ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OIi0liIIIoiOooLllLO0O0IoLLllIOlli ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OI0OLOILiOlOoolLIilooolollLLo0OOO ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( O0Il0L0lLloiIiliL0000o0oIOLLILool ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( Oo00IIIIoOIO0IL00llOoOioiollIOi00 ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OlIliOioiio0LLoLl00i0liioIOI00iIi ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OLOlLlooLIlL0IIiOilIiIooLloIioLOi ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOlOiiLoIooll0L00oIIIoOIililiillo ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( O0i000LoOoll00lolOOOOIO0Oio0LIO0o ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOiloioolOl0oLioOi0IoloOl0IlO0olL ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OlOlO00LLloOiOolOiOLOIiloLil0L0LI ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[18] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[18] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[18] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[18] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[18] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[18] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( Oo00OlooOo0io0OoIloiioLiOlL0llio0 ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OlIOlOillOlO0ol0iolIlLOiooOio0LOi ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OooOIi00Ii0liOollOoLioI0OiLiLiO0O ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OioolLOlII0IlolOIiLOliilL0oiiOoIo ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OoII0il0iLlL00iIo0I0OoloiiilLOLIo ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( Oi0Liloll0L00OiL0iLli0LO00iloIoLi ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OolIl0OOoiOlLioiloO0OolLOiIOolLLI ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOiiLLoL0llIoli0L0OOo0llL0oioiIlo ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[19] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[19] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[19] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[19] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[19] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[19] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OIl0oIiIIiLiIiLOiOOLOI0lOOOIIiIoo ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OOlO0o0i0Io0IOllLoIloiioiliOOlIII ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OO0llOooLooLoi0l0oIOOoilOolIoLLOo ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOIIlilOoOlIolLlILLioil0LL0oLlloo ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OOoooLL0l0llOLI0o0oO00LIoLO00LILO ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OoilLIlliloO0LoOL00IILioiolLIloi0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( Oll00iO0Ol0IOLloLLilo0OliIloIiLli ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OLllIIIO0oIlllOo00LILooILo0io0o00 ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OoI0LioOlolOLLL0iiIlOIooIlOoILLO0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OlOLIILoL0ll0oooOo0OIoLoOoiLIolol ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[20] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[20] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[20] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[20] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[20] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[20] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OOoOoILioOoIlIoLliOLOOi0io0IlLolo ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0oLiLiLlOlIIiLoLiLIiLL0l0oI0iIlO ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OIO0IioIOoIOIll0LOIlOOILoILoiilli ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLl0oiiIOL0ol00LIoo0IoolIollol0ii ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OiILIII00lOolOiililIOiIIloo0OlLlo ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O0lIi00lIl0iOlLilOloOIllllLLolooo ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OIl0iolIOLOlLOloIoLoIo0OooLi000lO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( Oiio0oo000ioIO0llioIoLILlIlIOOloL ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OoLOiILLiiloo0OOoOIOOooiLoiLoLiOI ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OIlLOILiLLo0ol0OLlI0IILilILLLlILO ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[21] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[21] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[21] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[21] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[21] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[21] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OiLllooo0Li0lioiolLi0ILIoLOliil0I ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0IL0iiIilolIlIiLIIIIOOiLOoOoloLL ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLoOLiILLLiIilOolo0Lil0iLLOOLILII ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O00liliooOOoiI0OlOOIIlO0o0IiOOolL ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OILLl0iillioLoOiiIiL0iliIOiO0oiio ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0I0LooLLiIO0illo0IliLLoioL0LlOLl ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OiioOooilOllI0oOoolilo0OLIlioo0II ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OIolOIIiLIloloOL0iIIO0il0li00ilOo ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OlOllIloiIIIIloliooOo0LoIil0o0oii ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OLILoOooIiil0oIIolILIlLIioL0i0Iio ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OIooL0lILLIloiOOLiI0ilOIli0LOL000 ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII Ol0IIiOloOLoOLlOiOo0LOoLIol0lOLOl ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[22] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[22] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[22] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[22] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[22] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[22] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0ILooiI0L00OoOoLlL0i0OooLOolooiO ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OlOlLO00i0Oiooo0lLollo0IILIlLO0OI ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOiOiIiiilililLoLlIOoIoiILilLoooI ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OIiolOOI00iliL0LolLOOOLOliiIlLlII ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0OoiooiIOLOllil0OLoLOlllL000LII0 ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OOl0i0OIIooLiI0IioL0LLILIloOlOllL ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OOOlLolILloIii0oollOil0lI0OOoOoo0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OOI0llLoO0IOO000OilllLLLI0i0Iilil ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOIOl00lliliioILLoiioolL0OLLoLo0i ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OII00III0LLIoI0LOloLoIo0IliiloOl0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[23] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[23] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[23] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[23] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[23] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[23] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OO0ooiOliiL0l0OoiiloO0oLIIIioII0L ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OLLliI0IiOiollllIOOLL0oL0IlllO0oI ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OO0O00OIoioOIOLi0IlILI0OlilooOIOo ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OlLo00LioOiOOOoliolIoLI0olOOlLoOI ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OLOL0OioiLOLoli0LOL00OOiO0iiOooll ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0oiOOLLiiillOliOOOllO0iO000OOoLI ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OIliOOilOillIo00oiOOLIOiLolIIooOl ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OIlOIiiliIlIOIlilliilOl0iILIOOOLO ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OIoll0OLiliiLlIililii0oiII0Ol00lO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( Ol0LliIIIIiOOILo0ooioLolOOOololIo ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OlollLLLoL0iiI0lool0OOOOIiOoolioL ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OllloLIILloiiiOill0lOLooilli0Llii ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OlI0LiIOLlllllL0OO0oLLII0ilILLoil ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OOiIlillllLOI0oOOoILlol0ILoIoOLil ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[24] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[24] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[24] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[24] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[24] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[24] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0iilOLolIOOlILi0iI0LLlLloiLO0L0O ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OLO00iLliol0LLIOOIIO0IiLIllO0IL0O ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OlLIiOlioIILOllO00lLiI0LiIlOloIiI ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OliiLi0oooOIo0L0lLoil0ooooi00I0ol ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OlIIloOL0iLIOLlOlLILlloiioloooILi ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OolOOLl0OlII0OiiloIloOO00IllliiLO ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OIliolloLooOi0OolOOi0ILOlIliLi0o0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OIILiOiLOO0IILI0llIOoooi0oLiiOioO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OLOILIii00lILOLoLIIlOiioll0ilOLii ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( O0IlliiI0l00iOLL0oLilIILo00lLIolo ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OII0Iill0IOLO000li0iL0iLoiIoOoliL ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OoIL0ll0llIOoI0IoIioiILILllLLOOOL ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OlILOIOO0IiOoioLi0LO0iolLIL0Ilol0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OOIiO0olO0OLlo0liIoiOioiIO00oOIiL ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[25] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[25] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[25] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[25] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[25] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[25] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OIILI00Loo0ooOiOL000Ilo00ool0I0oo ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( O0OII0Ili0ilol00OLOLoiOl0OlLo0liO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OlIli0IolOiL0LoliLloo0olllliIiO0O ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OO00il0IO0lLoiilIo0ioiOiOOlLloioL ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLoLOlol00olO0oo0LLlolI0OiLo0llLI ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OlIiO0llI0O0Li00OLIILiOLi00OiLioL ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OoL0LLOIlII0oLlloILillo0IOilOi0Il ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( O0o0OillO0LllooIiILLoilol0lii0liL ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OIO0L0iO0iLllOLILO0IoLliLolI00lLI ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OoOll0iOi0l0LiioLllOoliOoO00Lloil ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OiIoioILioOLl0io00oiOiO0liliOlOoO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OOI0I0II0oOOO0LiLoO0I00LloOllilIl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OlilOOiLOlI0Lll0oll0oLoI00OoIoOlI ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[26] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[26] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[26] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[26] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[26] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[26] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OLL0OiLILloil0IoOlLIIloLIiIlllLil ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OOooo0i0LloOLo00OIOIllLLiILOLLll0 ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OOL0lolilI0oIloIoIIILooo0lOLOlolI ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLolOilolLoloilIloOOiioIloiI0L0Lo ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( O0lIlL0lLL00000ioioloooIoiiiioi00 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( Oioo00O0OIloLlOil00lLiI0oIOOOoIio ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( O0oL00LOlilLooOoiil0oLL0iIillLlLL ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OOILlooOIliLloiliIOi00LIlLIoli000 ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OLOlILilLoI0liOiooL00OOlo0i0LiiiI ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( O0oOLILIoIlLOIIollLOoL00o0O00OiOo ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( O0OllOiIO00LliIOoLolo0loIiL0LiIlI ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOOOLL0II0ioIiIIoLOolIOLIoLooIill ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OOIioIlLoOL00lOliIIllL00illo0L00o ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OIOioIiIlLoiilIoLooIILIILIIIol00O ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[27] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[27] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[27] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[27] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[27] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[27] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OILI0LLillilOlllLil0ioLoIiliOoLLo ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OlLlL0ilOI0II0l0ILLIlIOLOoI0LiLIi ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( O0oIiILIIO0LOOil00IlIoLiIilO00ooI ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OiIL00IOiOiiI00oiio0lLOlooIiLiOio ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OOIIilloi0OiOoo0iI0LI0LI00oILiLio ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OLiloooloollOoil0LlolLolOILlO00Ol ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOLOIoliioI0oo0Ol0lOLiLLLoIioioi0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OlolLlliLo0O0l0lOOolL0ioI0O0Li00l ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[28] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[28] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[28] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[28] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[28] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[28] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( O0Ll0LoIi00OO0iolo0ILiolI0LOolooi ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OIO00IOolLoOoOL0ILI00i0olI0IiiOOo ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OIOio00oLLL0o00LO00LLoI0LlL0OILlO ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( O0illollo0oliIl0OolOoIlIILL0OIioO ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( O0Il00oIILloI0IL0LiOO0i0lIiIoolio ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OOilLILioilLIliOlOoilOOIolLLiLl0I ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OiOo0O0ooiioi00lloILL0oLLoILOiLiO ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OLLLI0L0OOoiLoIoLIOOIOLLoiloliIi0 ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( Oo0oI0oLOLlloloiiLIIol0LilOlOIliI ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[29] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[29] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[29] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[29] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[29] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[29] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OoIloII0oLiOLOLIllOL0iOoooOliOIii ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( Ool0o0OoOlOiL00i00O0iloIO0Lo00oOI ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLololIl0LoiLooLIloiooLli0LOOLLli ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OILllI0lillIoilOIoooOll0LII00I0l0 ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OLiILL00lIlOliLloi0OOl00LlIl0Loli ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OilIl00OOIloIli0LIIii00LIIlILiL0L ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OoOoIOoI0LILoIlIliLIioOooOOOIOoli ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OI00OLIIi0LioLLLLllooOiOl0iolOO0I ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OLIIl0o0liIOIooiOII0liO0oLllOI0oO ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OlOiOoL0i0i0L00OL00l00OOoL0OLILol ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OlLILiOolLl0ioiLiLlILiILLlIOllloI ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OiiILoLLoiliOOiOLOLiO0ioOIll0Oooo ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[30] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[30] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[30] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[30] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[30] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[30] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OIlOi0LL0LOLOLLL0LIIio0LLliiIoilo ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OIllOIIOiOol000OoLIL0lLl0L00iIIIL ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OlLiolooLilLlLiil0l0iiO0IOILool00 ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OIoolOll00LlI00l0oIOLLIOI0I0LIILo ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ) );
 OIIOlIO0ooOLLoll0il0IlOloL0oOIlII OOlO0LooL0ooliolL0i0i0iiLliOOl00I ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ( OoiLlL0oiiIloLOoloIL0oLii00IIIoII ) , .OoOi0O0oOoL0looLo0IoOllOOILiLooLl (OoOi0O0oOoL0looLo0IoOllOOILiLooLl[31] ), .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ( Oo0LLillol0loLIo0iOl0oOLlIOlILoIO[31] ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OilOIloOO0LiLoIL0IIILoIi0Loilll0I[31] ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0[31] ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO ( O0I0oI0I000LllOOI0L0lOlIl000LIioO[31] ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[31] ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( 4'd0 ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( 16'd0 ) , .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ( 1'd1 ) , .OOooLlloIiioOOO0LLILl0liiillLILol ( OilOOiiLIo0ooi0OLoliio0iooIooil0o ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ( OIoiIlOo00oL0iL0o0iooollLlilLoIIo ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( O0lolLi0olIioIiIooOLLLlioIooLIill ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OolLO0OOloooOIOiiOilL0IiILL0iol0I ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OL0looio0Loioi0ill0olOo0o00ioOOII ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( Ol0LioliiiiOil0liLiOiolioOo0oioii ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OO0oIOllioLiLlLLlii0ilL0OlIliIilO ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OLOllOoI0IolOloolLolO0lIiolLiIILi ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOILLooOOlllIILoIiIioLIOI0LOiLiLI ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ) );
 OLIi0oO0OOIIOllOoo000loIOil0OLi0O OLIi0oO0OOIIOllOoo000loIOil0OLi0O ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI (OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI ) , .OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL (OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL ) , .Oo0OiL0Lll000LlioLiooLOLloiLiliii (Oo0OiL0Lll000LlioLiooLOLloiLiliii ) , .OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI (OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI ) , .OioiIooIlil0liIiOIi0lLLIllOioioli (OioiIooIlil0liIiOIi0lLLIllOioioli ) , .OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 (OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 ) , .OlLloLOlOi0iIiLIlOlLio000LLOLILli (OlLloLOlOi0iIiLIlOlLio000LLOLILli ) , .OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 (OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 ) , .OOlILOLoilIOloioiIoOLI0L0ooLO0Lll (OOlILOLoilIOloioiIoOLI0L0ooLO0Lll ) , .OolOlIOiIIoII0ll0IllLoOiIllIilOoO (OolOlIOiIIoII0ll0IllLoOiIllIilOoO ) , .OOIiiol0IOILiLloOLiLOIIlIIolooOIO (OOIiiol0IOILiLloOLiLOIIlIIolooOIO ) , .OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO (OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO ) , .OILili00ILILlO0LIoLlll0oliLio0liL (OILili00ILILlO0LIoLlll0oliLio0liL ) , .OoILoooiioLLiIIIoiIoiOIO0OllIlIlL (OoILoooiioLLiIIIoiIoiOIO0OllIlIlL ) , .OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO (OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO ) , .OIiiiIlLolLIoIioOoOolloi0L0loLoIL (OIiiiIlLolLIoIioOoOolloi0L0loLoIL ) , .OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO (OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO ) , .O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II (O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II ) , .OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO (OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO ) , .OOlO0o0i0Io0IOllLoIloiioiliOOlIII (OOlO0o0i0Io0IOllLoIloiioiliOOlIII ) , .OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I (OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I ) , .O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 (O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 ) , .OlOlLO00i0Oiooo0lLollo0IILIlLO0OI (OlOlLO00i0Oiooo0lLollo0IILIlLO0OI ) , .OLLliI0IiOiollllIOOLL0oL0IlllO0oI (OLLliI0IiOiollllIOOLL0oL0IlllO0oI ) , .OLO00iLliol0LLIOOIIO0IiLIllO0IL0O (OLO00iLliol0LLIOOIIO0IiLIllO0IL0O ) , .O0OII0Ili0ilol00OLOLoiOl0OlLo0liO (O0OII0Ili0ilol00OLOLoiOl0OlLo0liO ) , .OOL0lolilI0oIloIoIIILooo0lOLOlolI (OOL0lolilI0oIloIoIIILooo0lOLOlolI ) , .OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll (OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll ) , .OIO00IOolLoOoOL0ILI00i0olI0IiiOOo (OIO00IOolLoOoOL0ILI00i0olI0IiiOOo ) , .OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO (OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO ) , .OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 (OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 ) , .OIoiIlOo00oL0iL0o0iooollLlilLoIIo (OIoiIlOo00oL0iL0o0iooollLlilLoIIo ) , .Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ) , .O0oill0llILOilo0i0LIoOLIoolL0Il0o (O0oill0llILOilo0i0LIoOLIoolL0Il0o ) , .OlliILlLOilOl0LO0O0OilooiIIiOi0Ll (OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ) , .OOLoL0looIOoioIoOooIoLIiIiLiLoiOl (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) , .OIoIooIolOilIOlooOlOIIOoilLioOIIO (OIoIooIolOilIOlooOlOIIOoilLioOIIO ) , .OiL0LolLLIOlliloII00llOil0oIlOiIo (OiL0LolLLIOlliloII00llOil0oIlOiIo ) , .O0llIOIliLOO0iiOoO0OO0lIOloLoII0I (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ) , .OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL ) , .OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo (OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ) , .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl ) , .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol ) , .O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo (O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ) , .OILIloOoilLIL00IIOoOilLOO0L0iiIOO (OILIloOoilLIL00IIOoOilLOO0L0iiIOO), .O0oLLi0Ill00l0lioiLioiooIllloIiIl (O0oLLi0Ill00l0lioiLioiooIllloIiIl), .OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 (OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ) , .O0Loo0iiI0OlLOlOIiILOooOOlIoioOli (O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ) , .OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI (OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ) , .OOiiILlloiOoI0OlilIOoiiLOOLol0IoI (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ) , .Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l (Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ) , .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI (OOLOoolOi0LIo0olO0loLllIlllIiiIiI ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI (OOOLiLOilooIi0Iio00ilILoLIILOoOoI ) , .OLLOooI0ILL00ILloiliILLLiioooLliI (OLLOooI0ILL00ILloiliILLLiioooLliI ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI (OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI (O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ) , .OilOOioILlOIIOL0iioIOIi0oloooOoLl (OilOOioILlOIIOL0iioIOIi0oloooOoLl ) , .OI00OiLolooiIIiiILoIliO0O0loolIlI (OI00OiLolooiIIiiILoIliO0O0loolIlI ) , .OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo (OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ) , .OoI0IoiILOOLILioiioIOoOLioiiOlIio (OoI0IoiILOOLILioiioIOoOLioiiOlIio ) , .OIIOLLOIlOlLoi0oiOioLilOiioiiliLO (OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ) , .O0OlOIIOOIOIioo00liool0iIiI0I0Lll (O0OlOIIOOIOIioo00liool0iIiI0I0Lll ) , .O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii (O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii ) , .OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l (OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l ) , .OIiOIl0O0OLllloOl0oOoLoIllIL0illO (OIiOIl0O0OLllloOl0oOoLoIllIL0illO ) , .Oi0loi0OllIlIoI0ILloIllILIO0IIo0I (Oi0loi0OllIlIoI0ILloIllILIO0IIo0I ) , .OoLOIol0OLIIiloO0oLoiliOl0LilIolI (OoLOIol0OLIIiloO0oLoiliOl0LilIolI ) , .OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i (OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i ) , .OOloOOOOiILOioIlIOO0oILilOLLL00OO (OOloOOOOiILOioIlIOO0oILilOLLL00OO ) , .OOIlIOO0IL0OoLli0IoliIioOOlIILlii (OOIlIOO0IL0OoLli0IoliIioOOlIILlii ) , .OioOlll0OooLLL0IIIIIli0ollooo0L0L (OioOlll0OooLLL0IIIIIli0ollooo0L0L ) , .OooOLOOliIlIOlio00OO0oloLoOi0lliO (OooOLOOliIlIOlio00OO0oloLoOi0lliO ) , .OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI (OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ) , .O0I0oI0I000LllOOI0L0lOlIl000LIioO (O0I0oI0I000LllOOI0L0lOlIl000LIioO ) , .OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO (OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO ) , .OLlOiiLlLoolliOiO0i0lOloio0L0oL00 (OLlOiiLlLoolliOiO0i0lOloio0L0oL00 ) , .OilOI0i0lloo0Lll000I0OIoIOI0lioiO (OilOI0i0lloo0Lll000I0OIoIOI0lioiO ) , .OlooiiLooL0L00oIIiioLloiIolOoOlLo (OlooiiLooL0L00oIIiioLloiIolOoOlLo ) , .OLo0LOlILllLILOIiiiL0LIlLIoLlO0II (OLo0LOlILllLILOIiiiL0LIlLIoLlO0II ) , .OiiOioOIO00LOOLilooiooo0olO0illo0 (OiiOioOIO00LOOLilooiooo0olO0illo0 ) , .OLl0LoLoii00oiOOoilollii000iIOlOI (OLl0LoLoii00oiOOoilollii000iIOlOI ) , .OLlil0000Oiil0IOOLiloIlliOoLLol0L (OLlil0000Oiil0IOOLiloIlliOoLLol0L ) , .OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI (OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI ) , .OO0OOILiO000LOILL0OllLi0l0oliLOo0 (OO0OOILiO000LOILL0OllLi0l0oliLOo0 ) , .OLiLllIIIlo0llILiLloLOoooOLOilI0l (OLiLllIIIlo0llILiLloLOoooOLOilI0l ) , .Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl (Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl ) , .OiL0IiiliiioOOLliLiiLILlIOloOLL0L (OiL0IiiliiioOOLliLiiLILlIOloOLL0L ) , .OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi (OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi ) , .OllLOLiIilI0oili000OiLilLioIOoIl0 (OllLOLiIilI0oili000OiLilLioIOoIl0 ) , .OOooI0loOL0iiOIoOili0OOOLLiiIiLOl (OOooI0loOL0iiOIoOili0OOOLLiiIiLOl ) , .OLIIiIIIOILl0loi0lO0IiOoolLIloi00 (OLIIiIIIOILl0loi0lO0IiOoolLIloi00 ) , .OoOillIILLoLoOioLloli0OLILlIOOoLo (OoOillIILLoLoOioLloli0OLILlIOOoLo ) , .OlOlO00LLloOiOolOiOLOIiloLil0L0LI (OlOlO00LLloOiOolOiOLOIiloLil0L0LI ) , .OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO (OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO ) , .OlOLIILoL0ll0oooOo0OIoLoOoiLIolol (OlOLIILoL0ll0oooOo0OIoLoOoiLIolol ) , .OIlLOILiLLo0ol0OLlI0IILilILLLlILO (OIlLOILiLLo0ol0OLlI0IILilILLLlILO ) , .O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i (O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i ) , .Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL (Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL ) , .OOiIlillllLOI0oOOoILlol0ILoIoOLil (OOiIlillllLOI0oOOoILlol0ILoIoOLil ) , .OOIiO0olO0OLlo0liIoiOioiIO00oOIiL (OOIiO0olO0OLlo0liIoiOioiIO00oOIiL ) , .O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 (O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 ) , .OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l (OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l ) , .OlolLlliLo0O0l0lOOolL0ioI0O0Li00l (OlolLlliLo0O0l0lOOolL0ioI0O0Li00l ) , .Oo0oI0oLOLlloloiiLIIol0LilOlOIliI (Oo0oI0oLOLlloloiiLIIol0LilOlOIliI ) , .OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo (OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo ) , .OoiLlL0oiiIloLOoloIL0oLii00IIIoII (OoiLlL0oiiIloLOoloIL0oLii00IIIoII ) , .Oo0LLillol0loLIo0iOl0oOLlIOlILoIO (Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ) , .OO0liOO0iOOIioool0OoLliiiI0l0ilOo (OO0liOO0iOOIioool0OoLliiiI0l0ilOo ) , .OiIOLi00lOILlOOL0oLLloL0io0LoIoOL (OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ) );
 Oi0IlLoiOlilloiLOloioOOiio0IiI0Io Oi0IlLoiOlilloiLOloioOOiio0IiI0Io ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OloliIooiiLI0IIlOiL0LLlioILLllL0L ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OioILlIiO0000OoolooO00loIOIloLIoI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLOl0000OLooLIIo0lIOIOI0lILioolOl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OoIolLlOIIoIoi00lloLlIoI0lo0iILol ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOIIloOlOILliIOILOIOiIlooIOOIL0oO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( O0liLooiLliIoLOllliIlo0ILo0I0oOOl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0i00oOl00OoIIOIil0LLOi0looIOIL00 ) , .OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ( OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ) , .OoolLolOioLILoOIII00LIOli00LIlloi ( OoolLolOioLILoOIII00LIOli00LIlloi ) , .OOOooLlOLO0iOOOLi00oIiloILlooOLIO ( OOOooLlOLO0iOOOLi00oIiloILlooOLIO ) , .OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ( OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ) , .OioLioLloIiilLLoOlIoiLIO0IOoiLoll ( OioLioLloIiilLLoOlIoiLIO0IOoiLoll ) , .Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ( Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ) , .OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ( OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ) , .OIiO0OLioLiIOIIiLoiLooI00I0olI00O ( OIiO0OLioLiIOIIiLoiLooI00I0olI00O ) , .OOOo0I0LlloiIl0i0il0OLiOlooOOolil ( OOOo0I0LlloiIl0i0il0OLiOlooOOolil ) , .OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ( OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ) , .OLlOlii00IoIl00oIioIiIool0lLiOoLo ( OLlOlii00IoIl00oIioIiIool0lLiOoLo ) , .OIollo0oLlLiI0IILOO00illIILLIoo0o ( OIollo0oLlLiI0IILOO00illIILLIoo0o ) , .O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ( O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ) , .OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ( OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ) , .OLli0lIO0lOO0OooILllIi00Lol00oili ( OLli0lIO0lOO0OooILllIi00Lol00oili ) , .Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ( Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ) , .OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ( OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ) , .OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ( OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ) , .OOIolooo0Oi00io00lIiiOiiLIliliOio ( OOIolooo0Oi00io00lIiiOiiLIliliOio ) , .OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ( OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ) , .O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ( O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ) , .OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ( OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ) , .OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ( OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ) , .Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ( Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ) , .O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ( O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ) , .OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ( OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ) , .OoI00LooIIlIIlIOOLIoloilI0OoIILLi ( OoI00LooIIlIIlIOOLIoloilI0OoIILLi ) , .OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ( OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ) , .O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ( O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ) , .OOIoOIilLi0looLILloOOollIIIo0llLo ( OOIoOIilLi0looLILloOOollIIIo0llLo ) , .OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ( OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ) , .OOllI0oo0L0io0l0IoloioOii0oIioOi0 ( OOllI0oo0L0io0l0IoloioOii0oIioOi0 ) , .OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ( OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ) , .Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ( Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ) , .O0oLiillllLOiLilOoI000iOLoiL0L0LO ( O0oLiillllLOiLilOoI000iOLoiL0L0LO ) , .OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ( OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ) , .Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ( Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ) , .OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ( OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ) , .OI0ioOlloiIio0oiOloi0lioiILoollLl ( OI0ioOlloiIio0oiOloi0lioiILoollLl ) , .OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ( OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ) , .OlIloooO00OIL0L0iIili0iOOoiLI0oiI ( OlIloooO00OIL0L0iIili0iOOoiLI0oiI ) , .OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ( OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ) , .OolIilIL0iooOLllOLloloOIlLIiOoLo0 ( OolIilIL0iooOLllOLloloOIlLIiOoLo0 ) , .OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ( OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ) , .OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ( OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ) , .O0lIOiilLOiIOollILlioiiOOiiLOO00i ( O0lIOiilLOiIOollILlioiiOOiiLOO00i ) , .O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ( O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ) , .OIiLIoliOIilIl0O00Li00oIO0OlIiooo ( OIiLIoliOIilIl0O00Li00oIO0OlIiooo ) , .OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ( OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ) , .O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ( O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ) , .Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ( Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ) , .Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ( Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ) , .OOoL0lOOloLLOLOILLLOolliIll0oOOoO ( OOoL0lOOloLLOLOILLLOolliIll0oOOoO ) , .OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ( OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ) , .OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ( OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ) , .O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ( O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ) , .OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ( OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ) , .O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ( O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ) , .O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ( O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ) , .OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ( OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ) , .OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ( OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ) , .Ol000OloII0LlIII00IIOIlOiioOo0Iii ( Ol000OloII0LlIII00IIOIlOiioOo0Iii ) , .OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ( OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ) , .OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ( OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ) , .OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ( OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ) , .OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ( OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ) , .OLLli0LLl0LlILOoi000iLoiiOOOLooLI ( OLLli0LLl0LlILOoi000iLoiiOOOLooLI ) , .OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ( OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ) , .OoooIiooOl0i0oliO0lio0IOo0iIILLLi ( OoooIiooOl0i0oliO0lio0IOo0iIILLLi ) , .OoOlILlliliiOI0OLLoOOl0000iIo0IIo ( OoOlILlliliiOI0OLLoOOl0000iIo0IIo ) , .OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ( OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ) , .O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ( O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ) , .OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ( OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ) , .OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ( OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ) , .OLolLol0lLIIlIillI000oIlilLLloOii ( OLolLol0lLIIlIillI000oIlilLLloOii ) , .OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ( OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ) , .OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ( OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ) , .OO0O0oOlliIoIOlooIO0lOLolIilLllIO ( OO0O0oOlliIoIOlooIO0lOLolIilLllIO ) , .O00I0iOoILll0oILl0ILloii0LIIOOiIO ( O00I0iOoILll0oILl0ILloii0LIIOOiIO ) , .OlolloloolOo0o0LLLIl00Li0iiLl00ol ( OlolloloolOo0o0LLLIl00Li0iiLl00ol ) , .OIIli0ilooIlOLI0lLO0Oi0IilILOolii ( OIIli0ilooIlOLI0lLO0Oi0IilILOolii ) , .OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ( OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ) , .OoOOLol000OllOLI0LO0LO0LoIliO0iiL ( OoOOLol000OllOLI0LO0LO0LoIliO0iiL ) , .OoIooi0LILolioIilliiol0I0iLoioIoi ( OoIooi0LILolioIilliiol0I0iLoioIoi ) , .OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ( OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ) , .OLlLoL0lO0oOIOolIIoiILIO0oOilooll ( OLlLoL0lO0oOIOolIIoiILIO0oOilooll ) , .O0iI0Lil0liLOLiILLOoilII0LII0iolO ( O0iI0Lil0liLOLiILLOoilII0LII0iolO ) , .OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ( OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ) , .OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ( OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ) , .O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ( O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ) , .OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ( OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ) , .OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ( OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ) , .OLLloO00IliLiLLlLloLloO0liOoIIOOI ( OLLloO00IliLiLLlLloLloO0liOoIIOOI ) , .OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ( OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ) , .OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ( OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ) , .OO00IIiOlOioiOLIiIloilLII0lLL0OOi ( OO00IIiOlOioiOLIiIloilLII0lLL0OOi ) , .OOLIlLlLIloIOoooilolooLloIi0OiiIi ( OOLIlLlLIloIOoooilolooLloIi0OiiIi ) , .OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ( OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ) , .OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ( OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ) , .OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ( OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ) , .OILolilliOIlLILOoioLii0iI0lII0oil ( OILolilliOIlLILOoioLii0iI0lII0oil ) , .OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ( OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ) , .OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ( OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ) , .O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ( O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ) , .OoLLliL00LLoooll00ooiLolOliOO0lLI ( OoLLliL00LLoooll00ooiLolOliOO0lLI ) , .OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ( OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ) , .O00loOoIIlII0OOo0lio00iOOOolLiIiO ( O00loOoIIlII0OOo0lio00iOOOolLiIiO ) , .OiiOIoolI0LioIo0IlL0lOllILIOOiIio ( OiiOIoolI0LioIo0IlL0lOllILIOOiIio ) , .OoIooolIllLIIolLII0IiLLiiOlOOIIOO ( OoIooolIllLIIolLII0IiLLiiOlOOIIOO ) , .OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ( OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ) , .OLL0i00LllLlio0oLOLooIL0ilLLllil0 ( OLL0i00LllLlio0oLOLooIL0ilLLllil0 ) , .OOiOiOIIoOii0oOLlI0OliIi0liioLLII ( OOiOiOIIoOii0oOLlI0OliIi0liioLLII ) , .OlOl0iOIioolOiill0OLOloOoLiIlllol ( OlOl0iOIioolOiill0OLOloOoLiIlllol ) , .OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ( OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ) , .OloILiOiLoIOOl0IoloOlI00Oollol0lL ( OloILiOiLoIOOl0IoloOlI00Oollol0lL ) , .OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ( OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ) , .OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ( OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ) , .OOIilioOiLLoOIL0iLoILiLLliiio0LOl ( OOIilioOiLLoOIL0iLoILiLLliiio0LOl ) , .O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ( O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ) , .Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ( Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ) , .O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ( O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ) , .O0li0llLIi0oIo0IilLLooLILolLIOOoo ( O0li0llLIi0oIo0IilLLooLILolLIOOoo ) , .OioIOIo0IllIo0OILLlli0LOOl00lioII ( OioIOIo0IllIo0OILLlli0LOOl00lioII ) , .OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ( OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ) , .OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ( OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ) , .Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ( Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ) , .OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ( OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ) , .OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ( OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ) , .O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ( O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ) , .OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ( OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ) , .OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ( OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ) , .O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ( O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ) , .OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ( OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ) , .OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ( OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ) , .OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ( OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ) , .OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ( OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ) , .Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ( Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ) , .O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ( O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ) , .OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ( OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ) , .O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ( O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ) , .O0il0OIIioo0IoL0OI0llOiLiLioill0i ( O0il0OIIioo0IoL0OI0llOiLiLioill0i ) , .O0lioOi00lO0IL00IoLLILolIlli00LiI ( O0lioOi00lO0IL00IoLLILolIlli00LiI ) , .OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ( OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ) , .OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ( OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ) , .OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ( OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ) , .OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ( OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ) , .OioOlIooLl0IL0LiioIlILIolO0o0ii0l ( OioOlIooLl0IL0LiioIlILIolO0o0ii0l ) , .OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ( OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ) , .OI0ILilL0olIiOoL0lOiiooolOOllIIIL ( OI0ILilL0olIiOoL0lOiiooolOOllIIIL ) , .O0000LloLiliiLOoIi0iLiLli0iloOOLI ( O0000LloLiliiLOoIi0iLiLli0iloOOLI ) , .OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ( OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ) , .OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ( OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ) , .OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ( OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ) , .OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ( OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ) , .OIO0IIi0OIooOiLOIII0lLolililiOIll ( OIO0IIi0OIooOiLOIII0lLolililiOIll ) , .OioilLoll0OiiOooiLiIOiL0LiilILII0 ( OioilLoll0OiiOooiLiIOiL0LiilILII0 ) , .OLoli0Li0i0oO0olOOilIliIio0LOoIIO ( OLoli0Li0i0oO0olOOilIliIio0LOoIIO ) , .OLLOoOIo0oiL0IOOO0lill0iloILllIOO ( OLLOoOIo0oiL0IOOO0lill0iloILllIOO ) , .OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ( OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ) , .OIILOOOOIOl00OoIollioiiliIilolLLl ( OIILOOOOIOl00OoIollioiiliIilolLLl ) , .OiooooLLoI0OLilIIil0ilooLo0OIloLl ( OiooooLLoI0OLilIIil0ilooLo0OIloLl ) , .O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ( O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ) , .OiLiiLILIoLilioiLolliOl0LI00LLil0 ( OiLiiLILIoLilioiLolliOl0LI00LLil0 ) , .Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ( Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ) , .Oloo0IIooolliliLOLoLoL0oI0LOliLlL ( Oloo0IIooolliliLOLoLoL0oI0LOliLlL ) , .OIiIIlooOiolooLoI0iLi0loLiloiLOll ( OIiIIlooOiolooLoI0iLi0loLiloiLOll ) , .OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ( OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ) , .OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ( OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ) , .OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ( OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ) , .OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ( OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ) , .Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ( Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ) , .OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ( OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ) , .Ol0OLoIiI0OloLIlillLOloLioIIL0III ( Ol0OLoIiI0OloLIlillLOloLioIIL0III ) , .OiILooool0OiolIOIIlO0LiOliIiIL0Ii ( OiILooool0OiolIOIIlO0LiOliIiIL0Ii ) , .OlLiiOLII0io0OLOOiIiiO0IIililoolo ( OlLiiOLII0io0OLOOiIiiO0IIililoolo ) , .OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ( OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ) , .OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ( OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ) , .OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ( OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ) , .OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ( OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ) , .OLlolloLliiLO0IlIlLo0lIiiloL00OOL ( OLlolloLliiLO0IlIlLo0lIiiloL00OOL ) , .OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ( OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ) , .O00oIiiOLOoilolOol0OIIOII00lllOIo ( O00oIiiOLOoilolOol0OIIOII00lllOIo ) , .OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ( OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ) , .OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ( OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ) , .Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ( Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ) , .OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ( OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ) , .OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ( OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ) , .OLi0ooOo0OlIllLOILllLL00lL00Liii0 ( OLi0ooOo0OlIllLOILllLL00lL00Liii0 ) , .OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ( OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ) , .Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ( Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ) , .OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ( OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ) , .Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ( Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ) , .Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ( Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ) , .OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ( OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ) , .OOOLilOolI0LILLIoloIiO00OiIiLiiIo ( OOOLilOolI0LILLIoloIiO00OiIiLiiIo ) , .OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ( OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ) , .OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ( OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ) , .OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ( OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ) , .OlLi0LOI0LoLioI0loilIlo00iliILIoi ( OlLi0LOI0LoLioI0loilIlo00iliILIoi ) , .OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ( OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ) , .OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ( OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ) , .OiOoiILoiIiIIoll0loilLl00Ll00O0iL ( OiOoiILoiIiIIoll0loilLl00Ll00O0iL ) , .OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ( OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ) , .OIlLiI0I0l0olLllLI0LliOOlllliLL0i ( OIlLiI0I0l0olLllLI0LliOOlllliLL0i ) , .OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ( OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ) , .OO0OOoLL0O0OOOllioILi0liilLLloiLO ( OO0OOoLL0O0OOOllioILi0liilLLloiLO ) , .OlLlliliOioioOIoiLOIOiOoiiioIOLOO ( OlLlliliOioioOIoiLOIOiOoiiioIOLOO ) , .OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ( OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ) , .OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ( OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ) , .OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ( OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ) , .OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ( OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ) , .OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ( OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ) , .OliliILl0LLiioool00L00LoLLILio0lO ( OliliILl0LLiioool00L00LoLLILio0lO ) , .OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ( OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ) , .OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ( OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ) , .OLioIOLOILilililoO0ililOi0oiIoo0o ( OLioIOLOILilililoO0ililOi0oiIoo0o ) , .OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ( OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ) , .Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ( Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ) , .Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ( Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ) , .OioIoIoo0iIIlOilLlIoILioo0I0lo00o ( OioIoIoo0iIIlOilLlIoILioo0I0lo00o ) , .O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ( O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ) , .OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ( OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ) , .OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ( OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ) , .OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ( OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ) , .O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ( O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ) , .OoLiLLooILIo0iol0OIoliLi0iiioiIlI ( OoLiLLooILIo0iol0OIoliLi0iiioiIlI ) , .OI0ool0i0ollOOoloL00L0LlLIO0LIliI ( OI0ool0i0ollOOoloL00L0LlLIO0LIliI ) , .Oo0loliLllliloIiliOi0lILloLI0ILlO ( Oo0loliLllliloIiliOi0lILloLI0ILlO ) , .Ooi0OL0i0IioliooLiI00OoiL00looOIL ( Ooi0OL0i0IioliooLiI00OoiL00looOIL ) , .OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ( OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ) , .OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ( OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ) , .OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ( OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ) , .OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ( OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ) , .OoOLolo0o0IOilOOLI0OoioLilIliI0lO ( OoOLolo0o0IOilOOLI0OoioLilIliI0lO ) , .O0o0OiliollLIi0IiLilIiOlLOOOLO00i ( O0o0OiliollLIi0IiLilIiOlLOOOLO00i ) , .OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ( OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ) , .OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ( OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ) , .OOIILlIiIOiOIi0o0li0lolol0LIoOliI ( OOIILlIiIOiOIi0o0li0lolol0LIoOliI ) , .OOIlIio0iILll00lliIIioiIiOLlLLi00 ( OOIlIio0iILll00lliIIioiIiOLlLLi00 ) , .OlIollIiLi0IlLiolloLOOL000Oo0l0II ( OlIollIiLi0IlLiolloLOOL000Oo0l0II ) , .OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ( OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ) , .OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ( OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ) , .OiiooiLLOL0iiO0oILoOlLoololiIIo0o ( OiiooiLLOL0iiO0oILoOlLoololiIIo0o ) , .OL0Lio0lIililolilllOL0Li0lIi0I0LI ( OL0Lio0lIililolilllOL0Li0lIi0I0LI ) , .O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ( O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ) , .OolL0oo00LOo0LOoLiILllLo0loOoIiii ( OolL0oo00LOo0LOoLiILllLo0loOoIiii ) , .OIOIOlilIolIlLOLlLlll0IiOIiILiOol ( OIOIOlilIolIlLOLlLlll0IiOIiILiOol ) , .OiloLLIlO00Il0oo0io0Iilliiil0OolO ( OiloLLIlO00Il0oo0io0Iilliiil0OolO ) , .O0oOL0illOloooo0ioIiOLOooLILllLl0 ( O0oOL0illOloooo0ioIiOLOooLILllLl0 ) , .Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ( Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ) , .OlOL0OLLooilLiOliIOIOOlIio00Oiili ( OlOL0OLLooilLiOliIOIOOlIio00Oiili ) , .OO0oolOlI0iloil0ooIolIioiol00I00I ( OO0oolOlI0iloil0ooIolIioiol00I00I ) , .O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ( O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ) , .OLI00Il0O0lI0OoLI0oIloiOIiiILIill ( OLI00Il0O0lI0OoLI0oIloiOIiiILIill ) , .OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ( OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ) , .OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ( OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ) , .O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ( O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ) , .OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ( OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ) , .OOoLol0oioL0looOlO0io0oIillil0iI0 ( OOoLol0oioL0looOlO0io0oIillil0iI0 ) , .OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ( OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ) , .OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ( OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ) , .O0oilLoOiOiLLi0Li0lLOIooIiliILlii ( O0oilLoOiOiLLi0Li0lLOIooIiliILlii ) , .O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ( O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ) , .OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ( OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ) , .OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ( OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ) , .OLiILioillIololIOILoOLlI0LILLliIL ( OLiILioillIololIOILoOLlI0LILLliIL ) , .OoOOillllIiloIOIILO0lL0LIl0iOlIII ( OoOOillllIiloIOIILO0lL0LIl0iOlIII ) , .OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ( OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ) , .OLIoIliI0LI0liL0i0IIIiLloL000l0lO ( OLIoIliI0LI0liL0i0IIIiLloL000l0lO ) , .Oo00OloiOIoLi00Oo0ooiololoOoooLLO ( Oo00OloiOIoLi00Oo0ooiololoOoooLLO ) , .Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ( Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ) , .Ollil0L0OlO0loio0OLiLILo0OioO0iOO ( Ollil0L0OlO0loio0OLiLILo0OioO0iOO ) , .OLio000LoL0lOol0oIiLlILLIlOLLOIlO ( OLio000LoL0lOol0oIiLlILLIlOLLOIlO ) , .OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ( OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ) , .OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ( OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ) , .OILIi00LOILOoLIiLloLiLIolliOoooIo ( OILIi00LOILOoLIiLloLiLIolliOoooIo ) , .OioilI0Oo0oOil0lIioiILIOLLLOLLioO ( OioilI0Oo0oOil0lIioiILIOLLLOLLioO ) , .OI0L0iIOilOi0LlILL0l0liiiil0lOIii ( OI0L0iIOilOi0LlILL0l0liiiil0lOIii ) , .OlIIioIIlILoli0oIiIl0l0IlOlloooll ( OlIIioIIlILoli0oIiIl0l0IlOlloooll ) , .O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ( O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ) , .OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ( OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ) , .OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ( OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ) , .Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ( Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ) , .OIOO0oiiIiiOILOOioiiO00OIl0lilllO ( OIOO0oiiIiiOILOOioiiO00OIl0lilllO ) , .OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ( OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ) , .OO0iLILOLioOioLOoLIOlOlo0oOIollll ( OO0iLILOLioOioLOoLIOlOlo0oOIollll ) , .OI00OlLIOIiOOiIliIooII00LLLllLLOO ( OI00OlLIOIiOOiIliIooII00LLLllLLOO ) , .OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ( OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ) , .O0L0O0ioooOOiLLlLLOLiioooILolII0o ( O0L0O0ioooOOiLLlLLOLiioooILolII0o ) , .OoiiooOo00OI0O0loiolLOLioIOiI0LoI ( OoiiooOo00OI0O0loiolLOLioIOiI0LoI ) , .OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ( OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ) , .O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ( O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ) , .OIi0liIIIoiOooLllLO0O0IoLLllIOlli ( OIi0liIIIoiOooLllLO0O0IoLLllIOlli ) , .OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ( OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ) , .OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ( OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ) , .OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ( OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ) , .OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ( OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ) , .OI0OLOILiOlOoolLIilooolollLLo0OOO ( OI0OLOILiOlOoolLIilooolollLLo0OOO ) , .O0Il0L0lLloiIiliL0000o0oIOLLILool ( O0Il0L0lLloiIiliL0000o0oIOLLILool ) , .OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ( OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ) , .Oo00IIIIoOIO0IL00llOoOioiollIOi00 ( Oo00IIIIoOIO0IL00llOoOioiollIOi00 ) , .OlIliOioiio0LLoLl00i0liioIOI00iIi ( OlIliOioiio0LLoLl00i0liioIOI00iIi ) , .OLOlLlooLIlL0IIiOilIiIooLloIioLOi ( OLOlLlooLIlL0IIiOilIiIooLloIioLOi ) , .OOlOiiLoIooll0L00oIIIoOIililiillo ( OOlOiiLoIooll0L00oIIIoOIililiillo ) , .O0i000LoOoll00lolOOOOIO0Oio0LIO0o ( O0i000LoOoll00lolOOOOIO0Oio0LIO0o ) , .OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ( OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ) , .Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ( Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ) , .OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ( OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ) , .O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ( O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ) , .O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ( O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ) , .O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ( O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ) , .OooOIi00Ii0liOollOoLioI0OiLiLiO0O ( OooOIi00Ii0liOollOoLioI0OiLiLiO0O ) , .OioolLOlII0IlolOIiLOliilL0oiiOoIo ( OioolLOlII0IlolOIiLOliilL0oiiOoIo ) , .OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ( OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ) , .OoII0il0iLlL00iIo0I0OoloiiilLOLIo ( OoII0il0iLlL00iIo0I0OoloiiilLOLIo ) , .OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ( OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ) , .Oi0Liloll0L00OiL0iLli0LO00iloIoLi ( Oi0Liloll0L00OiL0iLli0LO00iloIoLi ) , .OolIl0OOoiOlLioiloO0OolLOiIOolLLI ( OolIl0OOoiOlLioiloO0OolLOiIOolLLI ) , .OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ( OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ) , .OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ( OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ) , .OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ( OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ) , .Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ( Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ) , .OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ( OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ) , .OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ( OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ) , .O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ( O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ) , .OO0llOooLooLoi0l0oIOOoilOolIoLLOo ( OO0llOooLooLoi0l0oIOOoilOolIoLLOo ) , .OOIIlilOoOlIolLlILLioil0LL0oLlloo ( OOIIlilOoOlIolLlILLioil0LL0oLlloo ) , .OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ( OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ) , .OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ( OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ) , .OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ( OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ) , .OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ( OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ) , .Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ( Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ) , .OOoooLL0l0llOLI0o0oO00LIoLO00LILO ( OOoooLL0l0llOLI0o0oO00LIoLO00LILO ) , .OoilLIlliloO0LoOL00IILioiolLIloi0 ( OoilLIlliloO0LoOL00IILioiolLIloi0 ) , .OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ( OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ) , .O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ( O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ) , .OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ( OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ) , .Oll00iO0Ol0IOLloLLilo0OliIloIiLli ( Oll00iO0Ol0IOLloLLilo0OliIloIiLli ) , .OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ( OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ) , .OLllIIIO0oIlllOo00LILooILo0io0o00 ( OLllIIIO0oIlllOo00LILooILo0io0o00 ) , .OIO0IioIOoIOIll0LOIlOOILoILoiilli ( OIO0IioIOoIOIll0LOIlOOILoILoiilli ) , .Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ( Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ) , .OLl0oiiIOL0ol00LIoo0IoolIollol0ii ( OLl0oiiIOL0ol00LIoo0IoolIollol0ii ) , .OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ( OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ) , .OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ( OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ) , .OiILIII00lOolOiililIOiIIloo0OlLlo ( OiILIII00lOolOiililIOiIIloo0OlLlo ) , .OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ( OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ) , .OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ( OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ) , .OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ( OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ) , .OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ( OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ) , .OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ( OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ) , .O0lIi00lIl0iOlLilOloOIllllLLolooo ( O0lIi00lIl0iOlLilOloOIllllLLolooo ) , .OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ( OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ) , .O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ( O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ) , .OIl0iolIOLOlLOloIoLoIo0OooLi000lO ( OIl0iolIOLOlLOloIoLoIo0OooLi000lO ) , .Oiio0oo000ioIO0llioIoLILlIlIOOloL ( Oiio0oo000ioIO0llioIoLILlIlIOOloL ) , .OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ( OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ) , .OLoOLiILLLiIilOolo0Lil0iLLOOLILII ( OLoOLiILLLiIilOolo0Lil0iLLOOLILII ) , .O00liliooOOoiI0OlOOIIlO0o0IiOOolL ( O00liliooOOoiI0OlOOIIlO0o0IiOOolL ) , .OILLl0iillioLoOiiIiL0iliIOiO0oiio ( OILLl0iillioLoOiiIiL0iliIOiO0oiio ) , .OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ( OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ) , .O0I0LooLLiIO0illo0IliLLoioL0LlOLl ( O0I0LooLLiIO0illo0IliLLoioL0LlOLl ) , .OiioOooilOllI0oOoolilo0OLIlioo0II ( OiioOooilOllI0oOoolilo0OLIlioo0II ) , .OIolOIIiLIloloOL0iIIO0il0li00ilOo ( OIolOIIiLIloloOL0iIIO0il0li00ilOo ) , .OlOllIloiIIIIloliooOo0LoIil0o0oii ( OlOllIloiIIIIloliooOo0LoIil0o0oii ) , .OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ( OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ) , .OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ( OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ) , .OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ( OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ) , .OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ( OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ) , .OLILoOooIiil0oIIolILIlLIioL0i0Iio ( OLILoOooIiil0oIIolILIlLIioL0i0Iio ) , .OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ( OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ) , .OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ( OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ) , .OIooL0lILLIloiOOLiI0ilOIli0LOL000 ( OIooL0lILLIloiOOLiI0ilOIli0LOL000 ) , .O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ( O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ) , .OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ( OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ) , .O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ( O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ) , .OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ( OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ) , .OOiOiIiiilililLoLlIOoIoiILilLoooI ( OOiOiIiiilililLoLlIOoIoiILilLoooI ) , .OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ( OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ) , .OIiolOOI00iliL0LolLOOOLOliiIlLlII ( OIiolOOI00iliL0LolLOOOLOliiIlLlII ) , .O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ( O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ) , .O0OoiooiIOLOllil0OLoLOlllL000LII0 ( O0OoiooiIOLOllil0OLoLOlllL000LII0 ) , .Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ( Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ) , .OOl0i0OIIooLiI0IioL0LLILIloOlOllL ( OOl0i0OIIooLiI0IioL0LLILIloOlOllL ) , .OOOlLolILloIii0oollOil0lI0OOoOoo0 ( OOOlLolILloIii0oollOil0lI0OOoOoo0 ) , .O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ( O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ) , .O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ( O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ) , .OOI0llLoO0IOO000OilllLLLI0i0Iilil ( OOI0llLoO0IOO000OilllLLLI0i0Iilil ) , .OOIOl00lliliioILLoiioolL0OLLoLo0i ( OOIOl00lliliioILLoiioolL0OLLoLo0i ) , .OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ( OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ) , .OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ( OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ) , .OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ( OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ) , .Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ( Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ) , .OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ( OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ) , .OO0O00OIoioOIOLi0IlILI0OlilooOIOo ( OO0O00OIoioOIOLi0IlILI0OlilooOIOo ) , .OlLo00LioOiOOOoliolIoLI0olOOlLoOI ( OlLo00LioOiOOOoliolIoLI0olOOlLoOI ) , .OLOL0OioiLOLoli0LOL00OOiO0iiOooll ( OLOL0OioiLOLoli0LOL00OOiO0iiOooll ) , .OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ( OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ) , .O0oiOOLLiiillOliOOOllO0iO000OOoLI ( O0oiOOLLiiillOliOOOllO0iO000OOoLI ) , .OIliOOilOillIo00oiOOLIOiLolIIooOl ( OIliOOilOillIo00oiOOLIOiLolIIooOl ) , .OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ( OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ) , .OIlOIiiliIlIOIlilliilOl0iILIOOOLO ( OIlOIiiliIlIOIlilliilOl0iILIOOOLO ) , .OIoll0OLiliiLlIililii0oiII0Ol00lO ( OIoll0OLiliiLlIililii0oiII0Ol00lO ) , .Ol0LliIIIIiOOILo0ooioLolOOOololIo ( Ol0LliIIIIiOOILo0ooioLolOOOololIo ) , .OlollLLLoL0iiI0lool0OOOOIiOoolioL ( OlollLLLoL0iiI0lool0OOOOIiOoolioL ) , .O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ( O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ) , .OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ( OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ) , .OllloLIILloiiiOill0lOLooilli0Llii ( OllloLIILloiiiOill0lOLooilli0Llii ) , .OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ( OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ) , .OlLIiOlioIILOllO00lLiI0LiIlOloIiI ( OlLIiOlioIILOllO00lLiI0LiIlOloIiI ) , .OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ( OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ) , .OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ( OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ) , .OliiLi0oooOIo0L0lLoil0ooooi00I0ol ( OliiLi0oooOIo0L0lLoil0ooooi00I0ol ) , .O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ( O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ) , .OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ( OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ) , .OlIIloOL0iLIOLlOlLILlloiioloooILi ( OlIIloOL0iLIOLlOlLILlloiioloooILi ) , .OolOOLl0OlII0OiiloIloOO00IllliiLO ( OolOOLl0OlII0OiiloIloOO00IllliiLO ) , .O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ( O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ) , .OIliolloLooOi0OolOOi0ILOlIliLi0o0 ( OIliolloLooOi0OolOOi0ILOlIliLi0o0 ) , .Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ( Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ) , .OIILiOiLOO0IILI0llIOoooi0oLiiOioO ( OIILiOiLOO0IILI0llIOoooi0oLiiOioO ) , .OLOILIii00lILOLoLIIlOiioll0ilOLii ( OLOILIii00lILOLoLIIlOiioll0ilOLii ) , .O0IlliiI0l00iOLL0oLilIILo00lLIolo ( O0IlliiI0l00iOLL0oLilIILo00lLIolo ) , .OII0Iill0IOLO000li0iL0iLoiIoOoliL ( OII0Iill0IOLO000li0iL0iLoiIoOoliL ) , .OoIL0ll0llIOoI0IoIioiILILllLLOOOL ( OoIL0ll0llIOoI0IoIioiILILllLLOOOL ) , .OlIli0IolOiL0LoliLloo0olllliIiO0O ( OlIli0IolOiL0LoliLloo0olllliIiO0O ) , .OO00il0IO0lLoiilIo0ioiOiOOlLloioL ( OO00il0IO0lLoiilIo0ioiOiOOlLloioL ) , .OLoLOlol00olO0oo0LLlolI0OiLo0llLI ( OLoLOlol00olO0oo0LLlolI0OiLo0llLI ) , .OlIiO0llI0O0Li00OLIILiOLi00OiLioL ( OlIiO0llI0O0Li00OLIILiOLi00OiLioL ) , .OoL0LLOIlII0oLlloILillo0IOilOi0Il ( OoL0LLOIlII0oLlloILillo0IOilOi0Il ) , .OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ( OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ) , .OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ( OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ) , .OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ( OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ) , .O0o0OillO0LllooIiILLoilol0lii0liL ( O0o0OillO0LllooIiILLoilol0lii0liL ) , .OIO0L0iO0iLllOLILO0IoLliLolI00lLI ( OIO0L0iO0iLllOLILO0IoLliLolI00lLI ) , .OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ( OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ) , .OoOll0iOi0l0LiioLllOoliOoO00Lloil ( OoOll0iOi0l0LiioLllOoliOoO00Lloil ) , .OiIoioILioOLl0io00oiOiO0liliOlOoO ( OiIoioILioOLl0io00oiOiO0liliOlOoO ) , .OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ( OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ) , .OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ( OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ) , .OOI0I0II0oOOO0LiLoO0I00LloOllilIl ( OOI0I0II0oOOO0LiLoO0I00LloOllilIl ) , .OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ( OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ) , .OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ( OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ) , .OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ( OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ) , .OLolOilolLoloilIloOOiioIloiI0L0Lo ( OLolOilolLoloilIloOOiioIloiI0L0Lo ) , .O0lIlL0lLL00000ioioloooIoiiiioi00 ( O0lIlL0lLL00000ioioloooIoiiiioi00 ) , .Oioo00O0OIloLlOil00lLiI0oIOOOoIio ( Oioo00O0OIloLlOil00lLiI0oIOOOoIio ) , .O0oL00LOlilLooOoiil0oLL0iIillLlLL ( O0oL00LOlilLooOoiil0oLL0iIillLlLL ) , .OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ( OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ) , .OOILlooOIliLloiliIOi00LIlLIoli000 ( OOILlooOIliLloiliIOi00LIlLIoli000 ) , .OLOlILilLoI0liOiooL00OOlo0i0LiiiI ( OLOlILilLoI0liOiooL00OOlo0i0LiiiI ) , .O0oOLILIoIlLOIIollLOoL00o0O00OiOo ( O0oOLILIoIlLOIIollLOoL00o0O00OiOo ) , .O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ( O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ) , .OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ( OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ) , .O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ( O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ) , .O0OllOiIO00LliIOoLolo0loIiL0LiIlI ( O0OllOiIO00LliIOoLolo0loIiL0LiIlI ) , .OOOOLL0II0ioIiIIoLOolIOLIoLooIill ( OOOOLL0II0ioIiIIoLOolIOLIoLooIill ) , .OOIioIlLoOL00lOliIIllL00illo0L00o ( OOIioIlLoOL00lOliIIllL00illo0L00o ) , .OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ( OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ) , .Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ( Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ) , .O0oIiILIIO0LOOil00IlIoLiIilO00ooI ( O0oIiILIIO0LOOil00IlIoLiIilO00ooI ) , .OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ( OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ) , .OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ( OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ) , .OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ( OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ) , .Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ( Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ) , .OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ( OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ) , .OiIL00IOiOiiI00oiio0lLOlooIiLiOio ( OiIL00IOiOiiI00oiio0lLOlooIiLiOio ) , .OOIIilloi0OiOoo0iI0LI0LI00oILiLio ( OOIIilloi0OiOoo0iI0LI0LI00oILiLio ) , .Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ( Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ) , .OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ( OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ) , .O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ( O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ) , .Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ( Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ) , .Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ( Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ) , .OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ( OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ) , .OLiloooloollOoil0LlolLolOILlO00Ol ( OLiloooloollOoil0LlolLolOILlO00Ol ) , .O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ( O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ) , .OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ( OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ) , .OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ( OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ) , .OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ( OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ) , .OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ( OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ) , .O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ( O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ) , .OIOio00oLLL0o00LO00LLoI0LlL0OILlO ( OIOio00oLLL0o00LO00LLoI0LlL0OILlO ) , .OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ( OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ) , .O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ( O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ) , .OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ( OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ) , .OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ( OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ) , .O0illollo0oliIl0OolOoIlIILL0OIioO ( O0illollo0oliIl0OolOoIlIILL0OIioO ) , .O0Il00oIILloI0IL0LiOO0i0lIiIoolio ( O0Il00oIILloI0IL0LiOO0i0lIiIoolio ) , .OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ( OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ) , .OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ( OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ) , .OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ( OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ) , .OOilLILioilLIliOlOoilOOIolLLiLl0I ( OOilLILioilLIliOlOoilOOIolLLiLl0I ) , .OiOo0O0ooiioi00lloILL0oLLoILOiLiO ( OiOo0O0ooiioi00lloILL0oLLoILOiLiO ) , .OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ( OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ) , .OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ( OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ) , .OLololIl0LoiLooLIloiooLli0LOOLLli ( OLololIl0LoiLooLIloiooLli0LOOLLli ) , .OILllI0lillIoilOIoooOll0LII00I0l0 ( OILllI0lillIoilOIoooOll0LII00I0l0 ) , .OLiILL00lIlOliLloi0OOl00LlIl0Loli ( OLiILL00lIlOliLloi0OOl00LlIl0Loli ) , .OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ( OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ) , .OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ( OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ) , .OilIl00OOIloIli0LIIii00LIIlILiL0L ( OilIl00OOIloIli0LIIii00LIIlILiL0L ) , .OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ( OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ) , .OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ( OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ) , .OoOoIOoI0LILoIlIliLIioOooOOOIOoli ( OoOoIOoI0LILoIlIliLIioOooOOOIOoli ) , .OI00OLIIi0LioLLLLllooOiOl0iolOO0I ( OI00OLIIi0LioLLLLllooOiOl0iolOO0I ) , .OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ( OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ) , .OLIIl0o0liIOIooiOII0liO0oLllOI0oO ( OLIIl0o0liIOIooiOII0liO0oLllOI0oO ) , .OlOiOoL0i0i0L00OL00l00OOoL0OLILol ( OlOiOoL0i0i0L00OL00l00OOoL0OLILol ) , .OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ( OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ) , .OlLILiOolLl0ioiLiLlILiILLlIOllloI ( OlLILiOolLl0ioiLiLlILiILLlIOllloI ) , .OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ( OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ) , .OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ( OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ) , .OIllOIIOiOol000OoLIL0lLl0L00iIIIL ( OIllOIIOiOol000OoLIL0lLl0L00iIIIL ) , .OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ( OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ) , .OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ( OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ) , .OlLiolooLilLlLiil0l0iiO0IOILool00 ( OlLiolooLilLlLiil0l0iiO0IOILool00 ) , .OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ( OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ) , .OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ( OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ) , .OIoolOll00LlI00l0oIOLLIOI0I0LIILo ( OIoolOll00LlI00l0oIOLLIOI0I0LIILo ) , .OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ( OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ) , .OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ( OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ) , .OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ( OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ) , .OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ( OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ) , .Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ( Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ) , .OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ( OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ) , .OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ( OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ) , .OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ( OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ) , .O0lolLi0olIioIiIooOLLLlioIooLIill ( O0lolLi0olIioIiIooOLLLlioIooLIill ) , .OolLO0OOloooOIOiiOilL0IiILL0iol0I ( OolLO0OOloooOIOiiOilL0IiILL0iol0I ) , .OL0looio0Loioi0ill0olOo0o00ioOOII ( OL0looio0Loioi0ill0olOo0o00ioOOII ) , .Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ( Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ) , .Ol0LioliiiiOil0liLiOiolioOo0oioii ( Ol0LioliiiiOil0liLiOiolioOo0oioii ) , .Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ( Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ) , .OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ( OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ) , .OO0oIOllioLiLlLLlii0ilL0OlIliIilO ( OO0oIOllioLiLlLLlii0ilL0OlIliIilO ) , .OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ( OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ) , .OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ( OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ) , .OLOllOoI0IolOloolLolO0lIiolLiIILi ( OLOllOoI0IolOloolLolO0lIiolLiIILi ) , .OOILLooOOlllIILoIiIioLIOI0LOiLiLI ( OOILLooOOlllIILoIiIioLIOI0LOiLiLI ) , .O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ( O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ) , .OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ( OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ) , .Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ( Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ) , .OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ( OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ) , .O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ( O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ) , .OLlLLIloIliiIloOLloolLoIlLoi0iIoO (OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi), .OL0O0lL0lIILiOLLil0LoIIIlILLO00ll (OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 ), .OlLlOiIi0OoLiIlI0OO0loo0o0lOo0oIi (Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL), .OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI (OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI) );
 endmodule
 module Oi0IlLoiOlilloiLOloioOOiio0IiI0Io ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI , OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 , OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol , OloliIooiiLI0IIlOiL0LLlioILLllL0L , O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO , OioILlIiO0000OoolooO00loIOIloLIoI , OLOl0000OLooLIIo0lIOIOI0lILioolOl , OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII , OoIolLlOIIoIoi00lloLlIoI0lo0iILol , OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI , OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo , OOIIloOlOILliIOILOIOiIlooIOOIL0oO , OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io , OiLOo0loOI00OL0Ooio0OIIlOLiooLOII , OlLilll0ilOLI0IIoO0li0l0OlO00oLIO , O0liLooiLliIoLOllliIlo0ILo0I0oOOl , O0i00oOl00OoIIOIil0LLOi0looIOIL00 , OlllLl0L0L0iO0lIloilOOo0iIIiOo00o , OOlOIlooi0LiIlLiilOL0LloiII0I0oLo , O0oLiillllLOiLilOoI000iOLoiL0L0LO , Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL , OoooIiooOl0i0oliO0lio0IOo0iIILLLi , OLlLoL0lO0oOIOolIIoiILIO0oOilooll , OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl , Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o , Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 , OLooLooiioOiOo00LLooO0OLoI0iLiLI0 , Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo , OLi0ooOo0OlIllLOILllLL00lL00Liii0 , OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I , OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o , OOIlIio0iILll00lliIIioiIiOLlLLi00 , OOiOLoILiiIiOLoOOOl0iOolLLloLLLil , OLio000LoL0lOol0oIiLlILLIlOLLOIlO , OoiiooOo00OI0O0loiolLOLioIOiI0LoI , Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl , OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I , OIO0IioIOoIOIll0LOIlOOILoILoiilli , OLoOLiILLLiIilOolo0Lil0iLLOOLILII , OOoLoi0LlLLLoIIllLLLIli0OI0LlliII , OiLl00LLioIio0iLiOiIOOOlLIlilOIOi , OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 , OlIli0IolOiL0LoliLloo0olllliIiO0O , OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 , Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 , OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO , OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 , OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo , O0lolLi0olIioIiIooOLLLlioIooLIill , OoolLolOioLILoOIII00LIOli00LIlloi , OOIolooo0Oi00io00lIiiOiiLIliliOio , OLLIiolLOOOliIoiIi0oLLiOllooIoiiI , OOoL0lOOloLLOLOILLLOolliIll0oOOoO , OoOlILlliliiOI0OLLoOOl0000iIo0IIo , O0iI0Lil0liLOLiILLOoilII0LII0iolO , O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 , O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI , O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 , OIO0IIi0OIooOiLOIII0lLolililiOIll , OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 , OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl , OO0OOoLL0O0OOOllioILi0liilLLloiLO , OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 , OlIollIiLi0IlLiolloLOOL000Oo0l0II , O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO , OOoIIOoIl0LIOllIO0L0oLoOIOoooiill , OiOIOlILOi0lIoOiIOIoOIllLILLiIliL , OO0LO0iliiL0Oi0OIIloILLOiO0LLloli , O00OiooIolIi0oIoIiiLlO0IiIO0ooLio , Oo0i0IlILOo0ooOiIlLOoiioll0LilllO , O00liliooOOoiI0OlOOIIlO0o0IiOOolL , O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI , Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO , OlLIiOlioIILOllO00lLiI0LiIlOloIiI , OO00il0IO0lLoiilIo0ioiOiOOlLloioL , OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl , O0oIiILIIO0LOOil00IlIoLiIilO00ooI , OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l , OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 , OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 , OolLO0OOloooOIOiiOilL0IiILL0iol0I , OOOooLlOLO0iOOOLi00oIiloILlooOLIO , OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI , Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi , OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO , OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO , OlL0ioloIOIoOLILilIIlIiLo0oIliOLI , OoLLliL00LLoooll00ooiLolOliOO0lLI , O0li0llLIi0oIo0IilLLooLILolLIOOoo , OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl , OioilLoll0OiiOooiLiIOiL0LiilILII0 , Ol0OLoIiI0OloLIlillLOloLioIIL0III , Oi0lll0000oiiLo0lOolIi0ooOiiI0lio , OlLlliliOioioOIoiLOIOiOoiiioIOLOO , OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 , OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO , OoIIiLoIL0llOo00oIi0oLi00oiill0Ll , OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili , O0IIL0iIliIIolLLiioLIILlIoI0o0IOI , O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO , OO0llOooLooLoi0l0oIOOoilOolIoLLOo , OLl0oiiIOL0ol00LIoo0IoolIollol0ii , OILLl0iillioLoOiiIiL0iliIOiO0oiio , OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 , OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 , OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I , OLoLOlol00olO0oo0LLlolI0OiLo0llLI , OLolOilolLoloilIloOOiioIloiI0L0Lo , OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi , OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o , OLololIl0LoiLooLIloiooLli0LOOLLli , OIllOIIOiOol000OoLIL0lLl0L00iIIIL , OL0looio0Loioi0ill0olOo0o00ioOOII , OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o , O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi , OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi , OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 , O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO , OLLIool0I0IooOOIoliL0Oo0iL0L0lOol , OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi , OioIOIo0IllIo0OILLlli0LOOl00lioII , O0l0lloOLloIiI0o0LIoi0LOllOIlO0io , OLoli0Li0i0oO0olOOilIliIio0LOoIIO , OiILooool0OiolIOIIlO0LiOliIiIL0Ii , OLIIoIiliIoiioIoLoI0LllolIIlO0LOi , OIlI0I0IooLOLIlLLLIlli0o0LLl0illI , O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 , OLLiIlIOlII00l00l0LoLLilL0l0OOOLo , OOoLol0oioL0looOlO0io0oIillil0iI0 , OILIi00LOILOoLIiLloLiLIolliOoooIo , OIi0liIIIoiOooLllLO0O0IoLLllIOlli , O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI , OOIIlilOoOlIolLlILLioil0LL0oLlloo , OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 , OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL , OOiOiIiiilililLoLlIOoIoiILilLoooI , OO0O00OIoioOIOLi0IlILI0OlilooOIOo , OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO , OlIiO0llI0O0Li00OLIILiOLi00OiLioL , O0lIlL0lLL00000ioioloooIoiiiioi00 , OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 , OioLlLLli0IiOllll0l0LiIoLiLLLOL0L , OILllI0lillIoilOIoooOll0LII00I0l0 , OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL , Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI , OioLioLloIiilLLoOlIoiLIO0IOoiLoll , OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo , OI0ioOlloiIio0oiOloi0lioiILoollLl , O0L0Ll0OOOO0O0oLloilIliooOLlILoIL , OiL0l0OlOOOLiOIliO0lII0OliliioOo0 , O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l , O00loOoIIlII0OOo0lio00iOOOolLiIiO , OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI , O0il0OIIioo0IoL0OI0llOiLiLioill0i , OLLOoOIo0oiL0IOOO0lill0iloILllIOO , OlLiiOLII0io0OLOOiIiiO0IIililoolo , Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO , OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 , OoLiLLooILIo0iol0OIoliLi0iiioiIlI , OiiooiLLOL0iiO0oILoOlLoololiIIo0o , OOlILLi0LIOoLiill0I0LOIOiOLoOO00I , OioilI0Oo0oOil0lIioiILIOLLLOLLioO , OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I , O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi , OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo , OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi , O0I0LooLLiIO0illo0IliLLoioL0LlOLl , OliI0i0iIOiOoiII0olii0OOO0LIOiLLi , OlLo00LioOiOOOoliolIoLI0olOOlLoOI , OliiLi0oooOIo0L0lLoil0ooooi00I0ol , OoL0LLOIlII0oLlloILillo0IOilOi0Il , Oioo00O0OIloLlOil00lLiI0oIOOOoIio , OIoOOO00OOolil0OIiIlllOOOo0Oil0oo , O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL , OLiILL00lIlOliLloi0OOl00LlIl0Loli , OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli , Ol0LioliiiiOil0liLiOiolioOo0oioii , Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi , OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi , OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO , OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL , OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI , OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 , OiiOIoolI0LioIo0IlL0lOllILIOOiIio , OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l , O0lioOi00lO0IL00IoLLILolIlli00LiI , OOiiIi0oILLIllilLLLOiIi0Ii0lii0II , OoiOoio0IOIoOio0olOLllllOIlLIoiL0 , Oi00i0oL0iIiLll0o0o0l0loi000ioOOL , OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo , OI0ool0i0ollOOoloL00L0LlLIO0LIliI , OL0Lio0lIililolilllOL0Li0lIi0I0LI , OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 , OI0L0iIOilOi0LlILL0l0liiiil0lOIii , OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL , OooOIi00Ii0liOollOoLioI0OiLiLiO0O , OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol , OiILIII00lOolOiililIOiIIloo0OlLlo , OiioOooilOllI0oOoolilo0OLIlioo0II , OIiolOOI00iliL0LolLOOOLOliiIlLlII , OLOL0OioiLOLoli0LOL00OOiO0iiOooll , O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO , OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo , O0oL00LOlilLooOoiil0oLL0iIillLlLL , Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl , OIOio00oLLL0o00LO00LLoI0LlL0OILlO , OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 , OlLiolooLilLlLiil0l0iiO0IOILool00 , Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i , OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 , Oo000ooL0O00L0illOlOLOO0oilOIi0Ll , OlIloooO00OIL0L0iIili0iOOoiLI0oiI , O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL , OLolLol0lLIIlIillI000oIlilLLloOii , OoIoIO0O0oOoilLlI000OIllIIoI0ioIl , OoIooolIllLIIolLII0IiLLiiOlOOIIOO , Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio , OI0i0lOolo0oOILo00ll0LIIOiOOlIoii , OIILOOOOIOl00OoIollioiiliIilolLLl , OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 , OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L , OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L , Oo0loliLllliloIiliOi0lILloLI0ILlO , O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io , O0oilLoOiOiLLi0Li0lLOIooIiliILlii , OlIIioIIlILoli0oIiIl0l0IlOlloooll , OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO , OioolLOlII0IlolOIiLOliilL0oiiOoIo , OLIoilIIoI0Ol0Oll0I0LloliiLlolIII , OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 , OIolOIIiLIloloOL0iIIO0il0li00ilOo , O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO , OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L , OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl , OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL , OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L , OIL0OiIiiiOLliIioloLo0lLILolLoLL0 , OILLLoLI0LiOLilloOiLOIlILI0Io0l0o , OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl , OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI , OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 , OIiO0OLioLiIOIIiLoiLooI00I0olI00O , O0Ol0i0loLlooOIiLoOlIilLolOlio0ll , OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I , O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi , OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo , OLLloO00IliLiLLlLloLloO0liOoIIOOI , OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi , OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI , OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L , OiooooLLoI0OLilIIil0ilooLo0OIloLl , OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO , OOOLilOolI0LILLIoloIiO00OiIiLiiIo , OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l , Ooi0OL0i0IioliooLiI00OoiL00looOIL , OolL0oo00LOo0LOoLiILllLo0loOoIiii , O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l , O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I , OllLlOiLLooiILOiiOOlLlL0LOII0LLOL , OilO0i0Lll00Iolo00lOOLiLiOiLO0lio , OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 , OLOl00iiILoiI00i0lOlLOi00IOLLlOIL , OlOllIloiIIIIloliooOo0LoIil0o0oii , O0OoiooiIOLOllil0OLoLOlllL000LII0 , O0oiOOLLiiillOliOOOllO0iO000OOoLI , OlIIloOL0iLIOLlOlLILlloiioloooILi , OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l , OOILlooOIliLloiliIOi00LIlLIoli000 , OiIL00IOiOiiI00oiio0lLOlooIiLiOio , O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo , OilIl00OOIloIli0LIIii00LIIlILiL0L , OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I , OO0oIOllioLiLlLLlii0ilL0OlIliIilO , OOOo0I0LlloiIl0i0il0OLiOlooOOolil , OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li , OolIilIL0iooOLllOLloloOIlLIiOoLo0 , OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO , OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 , OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl , OLL0i00LllLlio0oLOLooIL0ilLLllil0 , OLLLllOIlLOioiIIoOIOiLOILOioLlLLo , OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I , O0iooIILOi0llLIIoILoo0ilIIIlooLI0 , OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 , OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl , OliliILl0LLiioool00L00LoLLILio0lO , OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O , OIOIOlilIolIlLOLlLlll0IiOIiILiOol , OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo , OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 , OI0OLOILiOlOoolLIilooolollLLo0OOO , OoII0il0iLlL00iIo0I0OoloiiilLOLIo , Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l , OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl , OLIoLi0ioO0OLLl0LlIOillIoili0OIOI , Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i , OIliOOilOillIo00oiOOLIOiLolIIooOl , OolOOLl0OlII0OiiloIloOO00IllliiLO , O0o0OillO0LllooIiILLoilol0lii0liL , OLOlILilLoI0liOiooL00OOlo0i0LiiiI , OOIIilloi0OiOoo0iI0LI0LI00oILiLio , OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 , OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O , OIoolOll00LlI00l0oIOLLIOI0I0LIILo , OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 , OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o , OoI00LooIIlIIlIOOLIoloilI0OoIILLi , OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII , OL0OIiOoo0IllO0oloolIll0oOo0LlIIi , OO0O0oOlliIoIOlooIO0lOLolIilLllIO , OOIlLIiol0o00OlI0lLl0lILiIolL0iIi , OOiOiOIIoOii0oOLlI0OliIi0liioLLII , O0oiILoiiI0oOOoiillLOoiIilI0o0Ool , OI0O0lOIO0OOOOllIL00Ooi0I0llLlili , OiLiiLILIoLilioiLolliOl0LI00LLil0 , OLlolloLliiLO0IlIlLo0lIiiloL00OOL , OooLI0lioLIOiOOI00oLLOiLIOlO00ILi , OL0Oloi0OoLOiO00LLloIolIo0iiLLOII , OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo , OiloLLIlO00Il0oo0io0Iilliiil0OolO , OLI0iO0OLLO00l00LIlOLiiLlloILOLIl , OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I , O0Il0L0lLloiIiliL0000o0oIOLLILool , OiI0ILIIIiiLO0LOlOLliioLL0II0OooL , OOoooLL0l0llOLI0o0oO00LIoLO00LILO , OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl , OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 , OOl0i0OIIooLiI0IioL0LLILIloOlOllL , OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO , O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O , OIO0L0iO0iLllOLILO0IoLliLolI00lLI , O0oOLILIoIlLOIIollLOoL00o0O00OiOo , Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl , OoooO0olOolLIIOLIIl0L0ooLIOoOOioL , OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o , OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 , OLoOO0OOIooLoI0liLOLllIiIOIL0Olol , OLlOlii00IoIl00oIioIiIool0lLiOoLo , OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL , OL0LLioOOooILOL0LLLIilLl0oLLiIoiL , Ol000OloII0LlIII00IIOIlOiioOo0Iii , O00I0iOoILll0oILl0ILloii0LIIOOiIO , OO00IIiOlOioiOLIiIloilLII0lLL0OOi , OlOl0iOIioolOiill0OLOloOoLiIlllol , OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 , OioOlIooLl0IL0LiioIlILIolO0o0ii0l , Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 , OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO , OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol , OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII , OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 , O0oOL0illOloooo0ioIiOLOooLILllLl0 , OLiILioillIololIOILoOLlI0LILLliIL , Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 , OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 , Oi0Liloll0L00OiL0iLli0LO00iloIoLi , OoilLIlliloO0LoOL00IILioiolLIloi0 , OLIloIl0iIiooOIo0lLlO0L00LOIil0LO , OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO , OOOlLolILloIii0oollOil0lI0OOoOoo0 , OIlOIiiliIlIOIlilliilOl0iILIOOOLO , OIliolloLooOi0OolOOi0ILOlIliLi0o0 , OI00OOL0LLOOLLLiIooi0oL0iioOloL0O , O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L , OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 , O0illollo0oliIl0OolOoIlIILL0OIioO , OoOoIOoI0LILoIlIliLIioOooOOOIOoli , OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L , OLOllOoI0IolOloolLolO0lIiolLiIILi , OIollo0oLlLiI0IILOO00illIILLIoo0o , O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 , O0lIOiilLOiIOollILlioiiOOiiLOO00i , OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I , OlolloloolOo0o0LLLIl00Li0iiLl00ol , OOLIlLlLIloIOoooilolooLloIi0OiiIi , OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO , OlIoO0LIi0LOLoLLOoliioiIOolIl00OO , OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI , Oloo0IIooolliliLOLoLoL0oI0LOliLlL , O00oIiiOLOoilolOol0OIIOII00lllOIo , OlLi0LOI0LoLioI0loilIlo00iliILIoi , OLioIOLOILilililoO0ililOi0oiIoo0o , OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL , Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo , OoOOillllIiloIOIILO0lL0LIl0iOlIII , OIOO0oiiIiiOILOOioiiO00OIl0lilllO , Oo00IIIIoOIO0IL00llOoOioiollIOi00 , OolIl0OOoiOlLioiloO0OolLOiIOolLLI , OL00oOoLi0iLl00LILOOLOlooiiLOOoLo , O0lIi00lIl0iOlLilOloOIllllLLolooo , OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL , O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 , OIoll0OLiliiLlIililii0oiII0Ol00lO , Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi , OoOll0iOi0l0LiioLllOoliOoO00Lloil , OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 , O00o0iOOoOiLI0iiIOoIiIliLoIliIIll , O0Il00oIILloI0IL0LiOO0i0lIiIoolio , OI00OLIIi0LioLLLLllooOiOl0iolOO0I , OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO , OOILLooOOlllIILoIiIioLIOI0LOiLiLI , O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL , OOIoOIilLi0looLILloOOollIIIo0llLo , O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL , OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll , OIIli0ilooIlOLI0lLO0Oi0IilILOolii , OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO , OloILiOiLoIOOl0IoloOlI00Oollol0lL , O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L , OI0ILilL0olIiOoL0lOiiooolOOllIIIL , OIiIIlooOiolooLoI0iLi0loLiloiLOll , OO0ilOiiOiIooOlIiO0l00iOliILoOIIi , OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO , OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL , OoOLolo0o0IOilOOLI0OoioLilIliI0lO , OlOL0OLLooilLiOliIOIOOlIio00Oiili , OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi , OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO , OlIliOioiio0LLoLl00i0liioIOI00iIi , OOiiILOoLlI00LoOil0OiOoIlloIiOi0o , O0ioLLo0liLOOiOL0OoLiOool0lLI00oi , OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o , OLILoOooIiil0oIIolILIlLIioL0i0Iio , O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O , Ol0LliIIIIiOOILo0ooioLolOOOololIo , OIILiOiLOO0IILI0llIOoooi0oLiiOioO , OiIoioILioOLl0io00oiOiO0liliOlOoO , O0OOOLLL0oOLoillIiOLIiIoI00LioiLl , Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo , OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO , OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO , OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO , O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi , OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi , OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL , OIiLIoliOIilIl0O00Li00oIO0OlIiooo , OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I , OlOlIILOLLIll0lo0lO0IOliliOOiL0oI , OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO , OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI , OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl , O0000LloLiliiLOoIi0iLiLli0iloOOLI , OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl , OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI , OI00ilIioiLo0ioiiIi0O0IolOiOi00IO , Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll , O0o0OiliollLIi0IiLilIiOlLOOOLO00i , OO0oolOlI0iloil0ooIolIioiol00I00I , OLIoIliI0LI0liL0i0IIIiLloL000l0lO , OO0iLILOLioOioLOoLIOlOlo0oOIollll , OLOlLlooLIlL0IIiOilIiIooLloIioLOi , OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 , OoIlL0lI0iL0iiIoLii0lLLio00lIIOol , O0O0L0iLLIlOILiOLoIiLiliiIllIi0li , OOLIlOoI0oOlII0oIllLi0l00iOioLIOi , OOI0llLoO0IOO000OilllLLLI0i0Iilil , OlollLLLoL0iiI0lool0OOOOIiOoolioL , OLOILIii00lILOLoLIIlOiioll0ilOLii , OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol , O0OllOiIO00LliIOoLolo0loIiL0LiIlI , Ooo00lolOl0OIoLOIlIliL0oLooIolLiL , OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol , OLIIl0o0liIOIooiOII0liO0oLllOI0oO , Olo0llLLi0L0IiLooLi0IooLOol0iIiIO , OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O , OLli0lIO0lOO0OooILllIi00Lol00oili , OOllI0oo0L0io0l0IoloioOii0oIioOi0 , OIIli0o0iiLOoOlilIoLIooOIooIL0ilI , OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio , OoOOLol000OllOLI0LO0LO0LoIliO0iiL , OoLOolIOLlOIIlIiOioiIIOL0lioliOIi , OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI , OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo , OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil , OI0IOio0lIIOiLllLLLIoIoiIoiOLillO , Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI , OiOoiILoiIiIIoll0loilLl00Ll00O0iL , Oo0IoILIliiOo0oooOLOiIo00i0L00Iio , OOooiloOoOIIiOiiLlLlLlIOIOIlolIol , O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI , Oo00OloiOIoLi00Oo0ooiololoOoooLLO , OI00OlLIOIiOOiIliIooII00LLLllLLOO , OOlOiiLoIooll0L00oIIIoOIililiillo , OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 , Oll00iO0Ol0IOLloLLilo0OliIloIiLli , OIl0iolIOLOlLOloIoLoIo0OooLi000lO , OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI , OOIOl00lliliioILLoiioolL0OLLoLo0i , O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 , O0IlliiI0l00iOLL0oLilIILo00lLIolo , OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl , OOOOLL0II0ioIiIIoLOolIOLIoLooIill , OLLI0ilo0LiioOLloOLloiioiIoOiLl0O , OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO , OlOiOoL0i0i0L00OL00l00OOoL0OLILol , OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO , Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l , Ooii00l0ooOoIliILL0lLLLLLoILlIIoO , OILl0LOii0lOi0LlLIIoIL0LLOoli0oll , O0Io0oIliooLo0i0i0lL0IlILOloiiIlI , OLLli0LLl0LlILOoi000iLoiiOOOLooLI , OoIooi0LILolioIilliiol0I0iLoioIoi , OILolilliOIlLILOoioLii0iI0lII0oil , OOIilioOiLLoOIL0iLoILiLLliiio0LOl , OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l , OllioLi0iLLoIOlILoIL0oOO0OiIliOOi , OlOoOLLlO0LOilOiiOoiOi0o0lollolLl , OILoioOioIOL0lIOLoIlIOlolLiOLlIoo , OoI0i0iiiL0ililIOLiL0IioLIL0IooOo , OioIoIoo0iIIlOilLlIoILioo0I0lo00o , OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 , OLI00Il0O0lI0OoLI0oIloiOIiiILIill , Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL , OioOiiiOlioLLOllo0IiIOiOOli0oi0LI , O0i000LoOoll00lolOOOOIO0Oio0LIO0o , Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO , OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl , Oiio0oo000ioIO0llioIoLILlIlIOOloL , OIooL0lILLIloiOOLiI0ilOIli0LOL000 , OILlOiiL00II0oiOlOoOI0lI00I0oIIIi , OLoOiiL00iolo0LOliOll0I0ILIOL0iLI , OII0Iill0IOLO000li0iL0iLoiIoOoliL , OOI0I0II0oOOO0LiLoO0I00LloOllilIl , OOIioIlLoOL00lOliIIllL00illo0L00o , OLiloooloollOoil0LlolLolOILlO00Ol , OOilLILioilLIliOlOoilOOIolLLiLl0I , OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 , OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI , OIiLOlOll0ol0OOLIo0oOiIilII0Io00L , OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI , Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO , Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi , OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI , OloIioIl0OOlolI0LIiioiLoL0OL0iI0i , OLIIoil00iiOOl0oloiiooOiI0IlL00Ol , O0L0oo0LI0OiII0l00oioIIiiilLLIOIl , OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl , OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo , OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI , OOoo0oiIolLIlol0oll00LiolIOOIlLL0 , OIlLiI0I0l0olLllLI0LliOOlllliLL0i , O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o , OOIILlIiIOiOIi0o0li0lolol0LIoOliI , OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL , Ollil0L0OlO0loio0OLiLILo0OioO0iOO , O0L0O0ioooOOiLLlLLOLiioooILolII0o , OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl , OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 , OLllIIIO0oIlllOo00LILooILo0io0o00 , OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI , O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO , OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 , OllloLIILloiiiOill0lOLooilli0Llii , OoIL0ll0llIOoI0IoIioiILILllLLOOOL , OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll , OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL , O0oLLI0O0IlOllolLIioIIOll0iiiIlLL , OiOo0O0ooiioi00lloILL0oLLoILOiLiO , OlLILiOolLl0ioiLiLlILiILLlIOllloI , OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O , O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi , OLlLLIloIliiIloOLloolLoIlLoi0iIoO, OL0O0lL0lIILiOLLil0LoIIIlILLO00ll , OlLlOiIi0OoLiIlI0OO0loo0o0lOo0oIi, OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI );
 parameter Ol0OioIIloLIlOLO0I0LoL0lIliIILI00 = 4'd0 ;
 parameter OiiOIloL0LLL0lO0lioLlL0o0LlL0IIOI = 4'd1 ;
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 input [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 input [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 input [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 input [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 input [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 input [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 input [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 input [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 input [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 input [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 input [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 input [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 input [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 input [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 input [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 input O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 input [ 23: 0] OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ;
 input [ 23: 0] OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ;
 input [ 23: 0] O0oLiillllLOiLilOoI000iOLoiL0L0LO ;
 input [ 23: 0] Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ;
 input [ 23: 0] OoooIiooOl0i0oliO0lio0IOo0iIILLLi ;
 input [ 23: 0] OLlLoL0lO0oOIOolIIoiILIO0oOilooll ;
 input [ 23: 0] OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ;
 input [ 23: 0] Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ;
 input [ 23: 0] Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ;
 input [ 23: 0] OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ;
 input [ 23: 0] Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ;
 input [ 23: 0] OLi0ooOo0OlIllLOILllLL00lL00Liii0 ;
 input [ 23: 0] OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ;
 input [ 23: 0] OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ;
 input [ 23: 0] OOIlIio0iILll00lliIIioiIiOLlLLi00 ;
 input [ 23: 0] OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ;
 input [ 23: 0] OLio000LoL0lOol0oIiLlILLIlOLLOIlO ;
 input [ 23: 0] OoiiooOo00OI0O0loiolLOLioIOiI0LoI ;
 input [ 23: 0] Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ;
 input [ 23: 0] OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ;
 input [ 23: 0] OIO0IioIOoIOIll0LOIlOOILoILoiilli ;
 input [ 23: 0] OLoOLiILLLiIilOolo0Lil0iLLOOLILII ;
 input [ 23: 0] OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ;
 input [ 23: 0] OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ;
 input [ 23: 0] OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ;
 input [ 23: 0] OlIli0IolOiL0LoliLloo0olllliIiO0O ;
 input [ 23: 0] OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ;
 input [ 23: 0] Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ;
 input [ 23: 0] OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ;
 input [ 23: 0] OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ;
 input [ 23: 0] OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ;
 input [ 23: 0] O0lolLi0olIioIiIooOLLLlioIooLIill ;
 input [ 7: 0] OoolLolOioLILoOIII00LIOli00LIlloi ;
 input [ 7: 0] OOIolooo0Oi00io00lIiiOiiLIliliOio ;
 input [ 7: 0] OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ;
 input [ 7: 0] OOoL0lOOloLLOLOILLLOolliIll0oOOoO ;
 input [ 7: 0] OoOlILlliliiOI0OLLoOOl0000iIo0IIo ;
 input [ 7: 0] O0iI0Lil0liLOLiILLOoilII0LII0iolO ;
 input [ 7: 0] O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ;
 input [ 7: 0] O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ;
 input [ 7: 0] O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ;
 input [ 7: 0] OIO0IIi0OIooOiLOIII0lLolililiOIll ;
 input [ 7: 0] OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ;
 input [ 7: 0] OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ;
 input [ 7: 0] OO0OOoLL0O0OOOllioILi0liilLLloiLO ;
 input [ 7: 0] OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ;
 input [ 7: 0] OlIollIiLi0IlLiolloLOOL000Oo0l0II ;
 input [ 7: 0] O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ;
 input [ 7: 0] OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ;
 input [ 7: 0] OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ;
 input [ 7: 0] OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ;
 input [ 7: 0] O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ;
 input [ 7: 0] Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ;
 input [ 7: 0] O00liliooOOoiI0OlOOIIlO0o0IiOOolL ;
 input [ 7: 0] O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ;
 input [ 7: 0] Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ;
 input [ 7: 0] OlLIiOlioIILOllO00lLiI0LiIlOloIiI ;
 input [ 7: 0] OO00il0IO0lLoiilIo0ioiOiOOlLloioL ;
 input [ 7: 0] OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ;
 input [ 7: 0] O0oIiILIIO0LOOil00IlIoLiIilO00ooI ;
 input [ 7: 0] OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ;
 input [ 7: 0] OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ;
 input [ 7: 0] OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ;
 input [ 7: 0] OolLO0OOloooOIOiiOilL0IiILL0iol0I ;
 input [ 31: 0] OOOooLlOLO0iOOOLi00oIiloILlooOLIO ;
 input [ 31: 0] OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ;
 input [ 31: 0] Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ;
 input [ 31: 0] OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ;
 input [ 31: 0] OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ;
 input [ 31: 0] OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ;
 input [ 31: 0] OoLLliL00LLoooll00ooiLolOliOO0lLI ;
 input [ 31: 0] O0li0llLIi0oIo0IilLLooLILolLIOOoo ;
 input [ 31: 0] OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ;
 input [ 31: 0] OioilLoll0OiiOooiLiIOiL0LiilILII0 ;
 input [ 31: 0] Ol0OLoIiI0OloLIlillLOloLioIIL0III ;
 input [ 31: 0] Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ;
 input [ 31: 0] OlLlliliOioioOIoiLOIOiOoiiioIOLOO ;
 input [ 31: 0] OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ;
 input [ 31: 0] OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ;
 input [ 31: 0] OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ;
 input [ 31: 0] OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ;
 input [ 31: 0] O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ;
 input [ 31: 0] O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ;
 input [ 31: 0] OO0llOooLooLoi0l0oIOOoilOolIoLLOo ;
 input [ 31: 0] OLl0oiiIOL0ol00LIoo0IoolIollol0ii ;
 input [ 31: 0] OILLl0iillioLoOiiIiL0iliIOiO0oiio ;
 input [ 31: 0] OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ;
 input [ 31: 0] OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ;
 input [ 31: 0] OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ;
 input [ 31: 0] OLoLOlol00olO0oo0LLlolI0OiLo0llLI ;
 input [ 31: 0] OLolOilolLoloilIloOOiioIloiI0L0Lo ;
 input [ 31: 0] OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ;
 input [ 31: 0] OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ;
 input [ 31: 0] OLololIl0LoiLooLIloiooLli0LOOLLli ;
 input [ 31: 0] OIllOIIOiOol000OoLIL0lLl0L00iIIIL ;
 input [ 31: 0] OL0looio0Loioi0ill0olOo0o00ioOOII ;
 input [ 7: 0] OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ;
 input [ 7: 0] O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ;
 input [ 7: 0] OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ;
 input [ 7: 0] OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ;
 input [ 7: 0] O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ;
 input [ 7: 0] OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ;
 input [ 7: 0] OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ;
 input [ 7: 0] OioIOIo0IllIo0OILLlli0LOOl00lioII ;
 input [ 7: 0] O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ;
 input [ 7: 0] OLoli0Li0i0oO0olOOilIliIio0LOoIIO ;
 input [ 7: 0] OiILooool0OiolIOIIlO0LiOliIiIL0Ii ;
 input [ 7: 0] OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ;
 input [ 7: 0] OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ;
 input [ 7: 0] O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ;
 input [ 7: 0] OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ;
 input [ 7: 0] OOoLol0oioL0looOlO0io0oIillil0iI0 ;
 input [ 7: 0] OILIi00LOILOoLIiLloLiLIolliOoooIo ;
 input [ 7: 0] OIi0liIIIoiOooLllLO0O0IoLLllIOlli ;
 input [ 7: 0] O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ;
 input [ 7: 0] OOIIlilOoOlIolLlILLioil0LL0oLlloo ;
 input [ 7: 0] OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ;
 input [ 7: 0] OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ;
 input [ 7: 0] OOiOiIiiilililLoLlIOoIoiILilLoooI ;
 input [ 7: 0] OO0O00OIoioOIOLi0IlILI0OlilooOIOo ;
 input [ 7: 0] OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ;
 input [ 7: 0] OlIiO0llI0O0Li00OLIILiOLi00OiLioL ;
 input [ 7: 0] O0lIlL0lLL00000ioioloooIoiiiioi00 ;
 input [ 7: 0] OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ;
 input [ 7: 0] OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ;
 input [ 7: 0] OILllI0lillIoilOIoooOll0LII00I0l0 ;
 input [ 7: 0] OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ;
 input [ 7: 0] Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ;
 input [ 31: 0] OioLioLloIiilLLoOlIoiLIO0IOoiLoll ;
 input [ 31: 0] OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ;
 input [ 31: 0] OI0ioOlloiIio0oiOloi0lioiILoollLl ;
 input [ 31: 0] O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ;
 input [ 31: 0] OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ;
 input [ 31: 0] O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ;
 input [ 31: 0] O00loOoIIlII0OOo0lio00iOOOolLiIiO ;
 input [ 31: 0] OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ;
 input [ 31: 0] O0il0OIIioo0IoL0OI0llOiLiLioill0i ;
 input [ 31: 0] OLLOoOIo0oiL0IOOO0lill0iloILllIOO ;
 input [ 31: 0] OlLiiOLII0io0OLOOiIiiO0IIililoolo ;
 input [ 31: 0] Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ;
 input [ 31: 0] OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ;
 input [ 31: 0] OoLiLLooILIo0iol0OIoliLi0iiioiIlI ;
 input [ 31: 0] OiiooiLLOL0iiO0oILoOlLoololiIIo0o ;
 input [ 31: 0] OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ;
 input [ 31: 0] OioilI0Oo0oOil0lIioiILIOLLLOLLioO ;
 input [ 31: 0] OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ;
 input [ 31: 0] O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ;
 input [ 31: 0] OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ;
 input [ 31: 0] OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ;
 input [ 31: 0] O0I0LooLLiIO0illo0IliLLoioL0LlOLl ;
 input [ 31: 0] OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ;
 input [ 31: 0] OlLo00LioOiOOOoliolIoLI0olOOlLoOI ;
 input [ 31: 0] OliiLi0oooOIo0L0lLoil0ooooi00I0ol ;
 input [ 31: 0] OoL0LLOIlII0oLlloILillo0IOilOi0Il ;
 input [ 31: 0] Oioo00O0OIloLlOil00lLiI0oIOOOoIio ;
 input [ 31: 0] OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ;
 input [ 31: 0] O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ;
 input [ 31: 0] OLiILL00lIlOliLloi0OOl00LlIl0Loli ;
 input [ 31: 0] OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ;
 input [ 31: 0] Ol0LioliiiiOil0liLiOiolioOo0oioii ;
 input [175: 0] Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ;
 input [175: 0] OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ;
 input [175: 0] OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ;
 input [175: 0] OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ;
 input [175: 0] OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ;
 input [175: 0] OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ;
 input [175: 0] OiiOIoolI0LioIo0IlL0lOllILIOOiIio ;
 input [175: 0] OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ;
 input [175: 0] O0lioOi00lO0IL00IoLLILolIlli00LiI ;
 input [175: 0] OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ;
 input [175: 0] OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ;
 input [175: 0] Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ;
 input [175: 0] OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ;
 input [175: 0] OI0ool0i0ollOOoloL00L0LlLIO0LIliI ;
 input [175: 0] OL0Lio0lIililolilllOL0Li0lIi0I0LI ;
 input [175: 0] OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ;
 input [175: 0] OI0L0iIOilOi0LlILL0l0liiiil0lOIii ;
 input [175: 0] OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ;
 input [175: 0] OooOIi00Ii0liOollOoLioI0OiLiLiO0O ;
 input [175: 0] OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ;
 input [175: 0] OiILIII00lOolOiililIOiIIloo0OlLlo ;
 input [175: 0] OiioOooilOllI0oOoolilo0OLIlioo0II ;
 input [175: 0] OIiolOOI00iliL0LolLOOOLOliiIlLlII ;
 input [175: 0] OLOL0OioiLOLoli0LOL00OOiO0iiOooll ;
 input [175: 0] O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ;
 input [175: 0] OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ;
 input [175: 0] O0oL00LOlilLooOoiil0oLL0iIillLlLL ;
 input [175: 0] Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ;
 input [175: 0] OIOio00oLLL0o00LO00LLoI0LlL0OILlO ;
 input [175: 0] OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ;
 input [175: 0] OlLiolooLilLlLiil0l0iiO0IOILool00 ;
 input [175: 0] Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ;
 input [ 71: 0] OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ;
 input [ 71: 0] Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ;
 input [ 71: 0] OlIloooO00OIL0L0iIili0iOOoiLI0oiI ;
 input [ 71: 0] O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ;
 input [ 71: 0] OLolLol0lLIIlIillI000oIlilLLloOii ;
 input [ 71: 0] OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ;
 input [ 71: 0] OoIooolIllLIIolLII0IiLLiiOlOOIIOO ;
 input [ 71: 0] Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ;
 input [ 71: 0] OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ;
 input [ 71: 0] OIILOOOOIOl00OoIollioiiliIilolLLl ;
 input [ 71: 0] OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ;
 input [ 71: 0] OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ;
 input [ 71: 0] OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ;
 input [ 71: 0] Oo0loliLllliloIiliOi0lILloLI0ILlO ;
 input [ 71: 0] O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ;
 input [ 71: 0] O0oilLoOiOiLLi0Li0lLOIooIiliILlii ;
 input [ 71: 0] OlIIioIIlILoli0oIiIl0l0IlOlloooll ;
 input [ 71: 0] OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ;
 input [ 71: 0] OioolLOlII0IlolOIiLOliilL0oiiOoIo ;
 input [ 71: 0] OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ;
 input [ 71: 0] OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ;
 input [ 71: 0] OIolOIIiLIloloOL0iIIO0il0li00ilOo ;
 input [ 71: 0] O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ;
 input [ 71: 0] OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ;
 input [ 71: 0] OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ;
 input [ 71: 0] OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ;
 input [ 71: 0] OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ;
 input [ 71: 0] OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ;
 input [ 71: 0] OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ;
 input [ 71: 0] OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ;
 input [ 71: 0] OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ;
 input [ 71: 0] OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ;
 input [ 31: 0] OIiO0OLioLiIOIIiLoiLooI00I0olI00O ;
 input [ 31: 0] O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ;
 input [ 31: 0] OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ;
 input [ 31: 0] O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ;
 input [ 31: 0] OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ;
 input [ 31: 0] OLLloO00IliLiLLlLloLloO0liOoIIOOI ;
 input [ 31: 0] OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ;
 input [ 31: 0] OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ;
 input [ 31: 0] OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ;
 input [ 31: 0] OiooooLLoI0OLilIIil0ilooLo0OIloLl ;
 input [ 31: 0] OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ;
 input [ 31: 0] OOOLilOolI0LILLIoloIiO00OiIiLiiIo ;
 input [ 31: 0] OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ;
 input [ 31: 0] Ooi0OL0i0IioliooLiI00OoiL00looOIL ;
 input [ 31: 0] OolL0oo00LOo0LOoLiILllLo0loOoIiii ;
 input [ 31: 0] O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ;
 input [ 31: 0] O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ;
 input [ 31: 0] OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ;
 input [ 31: 0] OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ;
 input [ 31: 0] OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ;
 input [ 31: 0] OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ;
 input [ 31: 0] OlOllIloiIIIIloliooOo0LoIil0o0oii ;
 input [ 31: 0] O0OoiooiIOLOllil0OLoLOlllL000LII0 ;
 input [ 31: 0] O0oiOOLLiiillOliOOOllO0iO000OOoLI ;
 input [ 31: 0] OlIIloOL0iLIOLlOlLILlloiioloooILi ;
 input [ 31: 0] OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ;
 input [ 31: 0] OOILlooOIliLloiliIOi00LIlLIoli000 ;
 input [ 31: 0] OiIL00IOiOiiI00oiio0lLOlooIiLiOio ;
 input [ 31: 0] O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ;
 input [ 31: 0] OilIl00OOIloIli0LIIii00LIIlILiL0L ;
 input [ 31: 0] OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ;
 input [ 31: 0] OO0oIOllioLiLlLLlii0ilL0OlIliIilO ;
 input [ 63: 0] OOOo0I0LlloiIl0i0il0OLiOlooOOolil ;
 input [ 63: 0] OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ;
 input [ 63: 0] OolIilIL0iooOLllOLloloOIlLIiOoLo0 ;
 input [ 63: 0] OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ;
 input [ 63: 0] OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ;
 input [ 63: 0] OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ;
 input [ 63: 0] OLL0i00LllLlio0oLOLooIL0ilLLllil0 ;
 input [ 63: 0] OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ;
 input [ 63: 0] OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ;
 input [ 63: 0] O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ;
 input [ 63: 0] OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ;
 input [ 63: 0] OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ;
 input [ 63: 0] OliliILl0LLiioool00L00LoLLILio0lO ;
 input [ 63: 0] OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ;
 input [ 63: 0] OIOIOlilIolIlLOLlLlll0IiOIiILiOol ;
 input [ 63: 0] OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ;
 input [ 63: 0] OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ;
 input [ 63: 0] OI0OLOILiOlOoolLIilooolollLLo0OOO ;
 input [ 63: 0] OoII0il0iLlL00iIo0I0OoloiiilLOLIo ;
 input [ 63: 0] Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ;
 input [ 63: 0] OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ;
 input [ 63: 0] OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ;
 input [ 63: 0] Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ;
 input [ 63: 0] OIliOOilOillIo00oiOOLIOiLolIIooOl ;
 input [ 63: 0] OolOOLl0OlII0OiiloIloOO00IllliiLO ;
 input [ 63: 0] O0o0OillO0LllooIiILLoilol0lii0liL ;
 input [ 63: 0] OLOlILilLoI0liOiooL00OOlo0i0LiiiI ;
 input [ 63: 0] OOIIilloi0OiOoo0iI0LI0LI00oILiLio ;
 input [ 63: 0] OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ;
 input [ 63: 0] OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ;
 input [ 63: 0] OIoolOll00LlI00l0oIOLLIOI0I0LIILo ;
 input [ 63: 0] OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ;
 input [ 31: 0] OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ;
 input [ 31: 0] OoI00LooIIlIIlIOOLIoloilI0OoIILLi ;
 input [ 31: 0] OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ;
 input [ 31: 0] OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ;
 input [ 31: 0] OO0O0oOlliIoIOlooIO0lOLolIilLllIO ;
 input [ 31: 0] OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ;
 input [ 31: 0] OOiOiOIIoOii0oOLlI0OliIi0liioLLII ;
 input [ 31: 0] O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ;
 input [ 31: 0] OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ;
 input [ 31: 0] OiLiiLILIoLilioiLolliOl0LI00LLil0 ;
 input [ 31: 0] OLlolloLliiLO0IlIlLo0lIiiloL00OOL ;
 input [ 31: 0] OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ;
 input [ 31: 0] OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ;
 input [ 31: 0] OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ;
 input [ 31: 0] OiloLLIlO00Il0oo0io0Iilliiil0OolO ;
 input [ 31: 0] OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ;
 input [ 31: 0] OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ;
 input [ 31: 0] O0Il0L0lLloiIiliL0000o0oIOLLILool ;
 input [ 31: 0] OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ;
 input [ 31: 0] OOoooLL0l0llOLI0o0oO00LIoLO00LILO ;
 input [ 31: 0] OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ;
 input [ 31: 0] OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ;
 input [ 31: 0] OOl0i0OIIooLiI0IioL0LLILIloOlOllL ;
 input [ 31: 0] OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ;
 input [ 31: 0] O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ;
 input [ 31: 0] OIO0L0iO0iLllOLILO0IoLliLolI00lLI ;
 input [ 31: 0] O0oOLILIoIlLOIIollLOoL00o0O00OiOo ;
 input [ 31: 0] Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ;
 input [ 31: 0] OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ;
 input [ 31: 0] OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ;
 input [ 31: 0] OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ;
 input [ 31: 0] OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ;
 input [ 63: 0] OLlOlii00IoIl00oIioIiIool0lLiOoLo ;
 input [ 63: 0] OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ;
 input [ 63: 0] OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ;
 input [ 63: 0] Ol000OloII0LlIII00IIOIlOiioOo0Iii ;
 input [ 63: 0] O00I0iOoILll0oILl0ILloii0LIIOOiIO ;
 input [ 63: 0] OO00IIiOlOioiOLIiIloilLII0lLL0OOi ;
 input [ 63: 0] OlOl0iOIioolOiill0OLOloOoLiIlllol ;
 input [ 63: 0] OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ;
 input [ 63: 0] OioOlIooLl0IL0LiioIlILIolO0o0ii0l ;
 input [ 63: 0] Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ;
 input [ 63: 0] OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ;
 input [ 63: 0] OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ;
 input [ 63: 0] OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ;
 input [ 63: 0] OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ;
 input [ 63: 0] O0oOL0illOloooo0ioIiOLOooLILllLl0 ;
 input [ 63: 0] OLiILioillIololIOILoOLlI0LILLliIL ;
 input [ 63: 0] Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ;
 input [ 63: 0] OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ;
 input [ 63: 0] Oi0Liloll0L00OiL0iLli0LO00iloIoLi ;
 input [ 63: 0] OoilLIlliloO0LoOL00IILioiolLIloi0 ;
 input [ 63: 0] OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ;
 input [ 63: 0] OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ;
 input [ 63: 0] OOOlLolILloIii0oollOil0lI0OOoOoo0 ;
 input [ 63: 0] OIlOIiiliIlIOIlilliilOl0iILIOOOLO ;
 input [ 63: 0] OIliolloLooOi0OolOOi0ILOlIliLi0o0 ;
 input [ 63: 0] OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ;
 input [ 63: 0] O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ;
 input [ 63: 0] OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ;
 input [ 63: 0] O0illollo0oliIl0OolOoIlIILL0OIioO ;
 input [ 63: 0] OoOoIOoI0LILoIlIliLIioOooOOOIOoli ;
 input [ 63: 0] OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ;
 input [ 63: 0] OLOllOoI0IolOloolLolO0lIiolLiIILi ;
 input [ 63: 0] OIollo0oLlLiI0IILOO00illIILLIoo0o ;
 input [ 63: 0] O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ;
 input [ 63: 0] O0lIOiilLOiIOollILlioiiOOiiLOO00i ;
 input [ 63: 0] OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ;
 input [ 63: 0] OlolloloolOo0o0LLLIl00Li0iiLl00ol ;
 input [ 63: 0] OOLIlLlLIloIOoooilolooLloIi0OiiIi ;
 input [ 63: 0] OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ;
 input [ 63: 0] OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ;
 input [ 63: 0] OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ;
 input [ 63: 0] Oloo0IIooolliliLOLoLoL0oI0LOliLlL ;
 input [ 63: 0] O00oIiiOLOoilolOol0OIIOII00lllOIo ;
 input [ 63: 0] OlLi0LOI0LoLioI0loilIlo00iliILIoi ;
 input [ 63: 0] OLioIOLOILilililoO0ililOi0oiIoo0o ;
 input [ 63: 0] OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ;
 input [ 63: 0] Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ;
 input [ 63: 0] OoOOillllIiloIOIILO0lL0LIl0iOlIII ;
 input [ 63: 0] OIOO0oiiIiiOILOOioiiO00OIl0lilllO ;
 input [ 63: 0] Oo00IIIIoOIO0IL00llOoOioiollIOi00 ;
 input [ 63: 0] OolIl0OOoiOlLioiloO0OolLOiIOolLLI ;
 input [ 63: 0] OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ;
 input [ 63: 0] O0lIi00lIl0iOlLilOloOIllllLLolooo ;
 input [ 63: 0] OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ;
 input [ 63: 0] O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ;
 input [ 63: 0] OIoll0OLiliiLlIililii0oiII0Ol00lO ;
 input [ 63: 0] Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ;
 input [ 63: 0] OoOll0iOi0l0LiioLllOoliOoO00Lloil ;
 input [ 63: 0] OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ;
 input [ 63: 0] O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ;
 input [ 63: 0] O0Il00oIILloI0IL0LiOO0i0lIiIoolio ;
 input [ 63: 0] OI00OLIIi0LioLLLLllooOiOl0iolOO0I ;
 input [ 63: 0] OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ;
 input [ 63: 0] OOILLooOOlllIILoIiIioLIOI0LOiLiLI ;
 input [ 63: 0] O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ;
 input [ 63: 0] OOIoOIilLi0looLILloOOollIIIo0llLo ;
 input [ 63: 0] O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ;
 input [ 63: 0] OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ;
 input [ 63: 0] OIIli0ilooIlOLI0lLO0Oi0IilILOolii ;
 input [ 63: 0] OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ;
 input [ 63: 0] OloILiOiLoIOOl0IoloOlI00Oollol0lL ;
 input [ 63: 0] O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ;
 input [ 63: 0] OI0ILilL0olIiOoL0lOiiooolOOllIIIL ;
 input [ 63: 0] OIiIIlooOiolooLoI0iLi0loLiloiLOll ;
 input [ 63: 0] OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ;
 input [ 63: 0] OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ;
 input [ 63: 0] OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ;
 input [ 63: 0] OoOLolo0o0IOilOOLI0OoioLilIliI0lO ;
 input [ 63: 0] OlOL0OLLooilLiOliIOIOOlIio00Oiili ;
 input [ 63: 0] OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ;
 input [ 63: 0] OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ;
 input [ 63: 0] OlIliOioiio0LLoLl00i0liioIOI00iIi ;
 input [ 63: 0] OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ;
 input [ 63: 0] O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ;
 input [ 63: 0] OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ;
 input [ 63: 0] OLILoOooIiil0oIIolILIlLIioL0i0Iio ;
 input [ 63: 0] O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ;
 input [ 63: 0] Ol0LliIIIIiOOILo0ooioLolOOOololIo ;
 input [ 63: 0] OIILiOiLOO0IILI0llIOoooi0oLiiOioO ;
 input [ 63: 0] OiIoioILioOLl0io00oiOiO0liliOlOoO ;
 input [ 63: 0] O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ;
 input [ 63: 0] Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ;
 input [ 63: 0] OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ;
 input [ 63: 0] OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ;
 input [ 63: 0] OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ;
 input [ 63: 0] O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ;
 input [ 31: 0] OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ;
 input [ 31: 0] OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ;
 input [ 31: 0] OIiLIoliOIilIl0O00Li00oIO0OlIiooo ;
 input [ 31: 0] OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ;
 input [ 31: 0] OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ;
 input [ 31: 0] OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ;
 input [ 31: 0] OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ;
 input [ 31: 0] OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ;
 input [ 31: 0] O0000LloLiliiLOoIi0iLiLli0iloOOLI ;
 input [ 31: 0] OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ;
 input [ 31: 0] OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ;
 input [ 31: 0] OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ;
 input [ 31: 0] Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ;
 input [ 31: 0] O0o0OiliollLIi0IiLilIiOlLOOOLO00i ;
 input [ 31: 0] OO0oolOlI0iloil0ooIolIioiol00I00I ;
 input [ 31: 0] OLIoIliI0LI0liL0i0IIIiLloL000l0lO ;
 input [ 31: 0] OO0iLILOLioOioLOoLIOlOlo0oOIollll ;
 input [ 31: 0] OLOlLlooLIlL0IIiOilIiIooLloIioLOi ;
 input [ 31: 0] OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ;
 input [ 31: 0] OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ;
 input [ 31: 0] O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ;
 input [ 31: 0] OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ;
 input [ 31: 0] OOI0llLoO0IOO000OilllLLLI0i0Iilil ;
 input [ 31: 0] OlollLLLoL0iiI0lool0OOOOIiOoolioL ;
 input [ 31: 0] OLOILIii00lILOLoLIIlOiioll0ilOLii ;
 input [ 31: 0] OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ;
 input [ 31: 0] O0OllOiIO00LliIOoLolo0loIiL0LiIlI ;
 input [ 31: 0] Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ;
 input [ 31: 0] OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ;
 input [ 31: 0] OLIIl0o0liIOIooiOII0liO0oLllOI0oO ;
 input [ 31: 0] Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ;
 input [ 31: 0] OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ;
 input [ 63: 0] OLli0lIO0lOO0OooILllIi00Lol00oili ;
 input [ 63: 0] OOllI0oo0L0io0l0IoloioOii0oIioOi0 ;
 input [ 63: 0] OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ;
 input [ 63: 0] OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ;
 input [ 63: 0] OoOOLol000OllOLI0LO0LO0LoIliO0iiL ;
 input [ 63: 0] OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ;
 input [ 63: 0] OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ;
 input [ 63: 0] OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ;
 input [ 63: 0] OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ;
 input [ 63: 0] OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ;
 input [ 63: 0] Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ;
 input [ 63: 0] OiOoiILoiIiIIoll0loilLl00Ll00O0iL ;
 input [ 63: 0] Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ;
 input [ 63: 0] OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ;
 input [ 63: 0] O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ;
 input [ 63: 0] Oo00OloiOIoLi00Oo0ooiololoOoooLLO ;
 input [ 63: 0] OI00OlLIOIiOOiIliIooII00LLLllLLOO ;
 input [ 63: 0] OOlOiiLoIooll0L00oIIIoOIililiillo ;
 input [ 63: 0] OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ;
 input [ 63: 0] Oll00iO0Ol0IOLloLLilo0OliIloIiLli ;
 input [ 63: 0] OIl0iolIOLOlLOloIoLoIo0OooLi000lO ;
 input [ 63: 0] OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ;
 input [ 63: 0] OOIOl00lliliioILLoiioolL0OLLoLo0i ;
 input [ 63: 0] O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ;
 input [ 63: 0] O0IlliiI0l00iOLL0oLilIILo00lLIolo ;
 input [ 63: 0] OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ;
 input [ 63: 0] OOOOLL0II0ioIiIIoLOolIOLIoLooIill ;
 input [ 63: 0] OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ;
 input [ 63: 0] OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ;
 input [ 63: 0] OlOiOoL0i0i0L00OL00l00OOoL0OLILol ;
 input [ 63: 0] OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ;
 input [ 63: 0] Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ;
 input [ 31: 0] Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ;
 input [ 31: 0] OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ;
 input [ 31: 0] O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ;
 input [ 31: 0] OLLli0LLl0LlILOoi000iLoiiOOOLooLI ;
 input [ 31: 0] OoIooi0LILolioIilliiol0I0iLoioIoi ;
 input [ 31: 0] OILolilliOIlLILOoioLii0iI0lII0oil ;
 input [ 31: 0] OOIilioOiLLoOIL0iLoILiLLliiio0LOl ;
 input [ 31: 0] OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ;
 input [ 31: 0] OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ;
 input [ 31: 0] OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ;
 input [ 31: 0] OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ;
 input [ 31: 0] OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ;
 input [ 31: 0] OioIoIoo0iIIlOilLlIoILioo0I0lo00o ;
 input [ 31: 0] OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ;
 input [ 31: 0] OLI00Il0O0lI0OoLI0oIloiOIiiILIill ;
 input [ 31: 0] Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ;
 input [ 31: 0] OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ;
 input [ 31: 0] O0i000LoOoll00lolOOOOIO0Oio0LIO0o ;
 input [ 31: 0] Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ;
 input [ 31: 0] OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ;
 input [ 31: 0] Oiio0oo000ioIO0llioIoLILlIlIOOloL ;
 input [ 31: 0] OIooL0lILLIloiOOLiI0ilOIli0LOL000 ;
 input [ 31: 0] OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ;
 input [ 31: 0] OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ;
 input [ 31: 0] OII0Iill0IOLO000li0iL0iLoiIoOoliL ;
 input [ 31: 0] OOI0I0II0oOOO0LiLoO0I00LloOllilIl ;
 input [ 31: 0] OOIioIlLoOL00lOliIIllL00illo0L00o ;
 input [ 31: 0] OLiloooloollOoil0LlolLolOILlO00Ol ;
 input [ 31: 0] OOilLILioilLIliOlOoilOOIolLLiLl0I ;
 input [ 31: 0] OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ;
 input [ 31: 0] OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ;
 input [ 31: 0] OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ;
 input OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ;
 input Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ;
 input Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ;
 input OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ;
 input OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ;
 input OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ;
 input O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ;
 input OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ;
 input OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ;
 input OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ;
 input OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ;
 input OIlLiI0I0l0olLllLI0LliOOlllliLL0i ;
 input O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ;
 input OOIILlIiIOiOIi0o0li0lolol0LIoOliI ;
 input OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ;
 input Ollil0L0OlO0loio0OLiLILo0OioO0iOO ;
 input O0L0O0ioooOOiLLlLLOLiioooILolII0o ;
 input OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ;
 input OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ;
 input OLllIIIO0oIlllOo00LILooILo0io0o00 ;
 input OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ;
 input O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ;
 input OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ;
 input OllloLIILloiiiOill0lOLooilli0Llii ;
 input OoIL0ll0llIOoI0IoIioiILILllLLOOOL ;
 input OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ;
 input OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ;
 input O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ;
 input OiOo0O0ooiioi00lloILL0oLLoILOiLiO ;
 input OlLILiOolLl0ioiLiLlILiILLlIOllloI ;
 input OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ;
 input O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ;
 output OLlLLIloIliiIloOLloolLoIlLoi0iIoO;
 output reg [255:0] OL0O0lL0lIILiOLLil0LoIIIlILLO00ll ;
 output reg OlLlOiIi0OoLiIlI0OO0loo0o0lOo0oIi;
 input OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI;
 wire [255:0] OlolI00LoLoOILILoioLOL0lolLO0oiOo ;
 wire [255:0] OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL ;
 wire [255:0] O0000Lil0OoOOILlIlOlooioiIOloOioi ;
 wire [ 31:0] O00lOOl0oILIoiioLOOI0OoioILioLiiL ;
 wire O0iioiILo0ol0ollLilLl0lO0oI0ilOiL ;
 wire [255:0] OilO0OLOo0LllI00o0oOil00L0OloIOl0 ;
 wire [255:0] OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll ;
 wire OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l ;
 wire OILLiiO0o00OloIOOl0LlIOOlo00O0OOi ;
 wire [255:0] OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil ;
 wire [255:0] Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 ;
 wire OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl ;
 wire Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI ;
 OlLIO0oiil0ooIiOOioiLOI0oooilILoi OlLIO0oiil0ooIiOOioiLOI0oooilILoi ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi ) , .OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ( OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ) , .OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ( OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ) , .OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ( OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ) , .OloliIooiiLI0IIlOiL0LLlioILLllL0L ( OloliIooiiLI0IIlOiL0LLlioILLllL0L ) , .O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ( O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ) , .OioILlIiO0000OoolooO00loIOIloLIoI ( OioILlIiO0000OoolooO00loIOIloLIoI ) , .OLOl0000OLooLIIo0lIOIOI0lILioolOl ( OLOl0000OLooLIIo0lIOIOI0lILioolOl ) , .OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ( OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ) , .OoIolLlOIIoIoi00lloLlIoI0lo0iILol ( OoIolLlOIIoIoi00lloLlIoI0lo0iILol ) , .OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ( OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ) , .OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ( OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ) , .OOIIloOlOILliIOILOIOiIlooIOOIL0oO ( OOIIloOlOILliIOILOIOiIlooIOOIL0oO ) , .OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ( OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ) , .OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ( OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ) , .OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ( OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ) , .O0liLooiLliIoLOllliIlo0ILo0I0oOOl ( O0liLooiLliIoLOllliIlo0ILo0I0oOOl ) , .O0i00oOl00OoIIOIil0LLOi0looIOIL00 ( O0i00oOl00OoIIOIil0LLOi0looIOIL00 ) , .OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ( OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ) , .OoolLolOioLILoOIII00LIOli00LIlloi ( OoolLolOioLILoOIII00LIOli00LIlloi ) , .OOOooLlOLO0iOOOLi00oIiloILlooOLIO ( OOOooLlOLO0iOOOLi00oIiloILlooOLIO ) , .OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ( OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ) , .OioLioLloIiilLLoOlIoiLIO0IOoiLoll ( OioLioLloIiilLLoOlIoiLIO0IOoiLoll ) , .Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ( Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ) , .OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ( OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ) , .OIiO0OLioLiIOIIiLoiLooI00I0olI00O ( OIiO0OLioLiIOIIiLoiLooI00I0olI00O ) , .OOOo0I0LlloiIl0i0il0OLiOlooOOolil ( OOOo0I0LlloiIl0i0il0OLiOlooOOolil ) , .OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ( OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ) , .OLlOlii00IoIl00oIioIiIool0lLiOoLo ( OLlOlii00IoIl00oIioIiIool0lLiOoLo ) , .OIollo0oLlLiI0IILOO00illIILLIoo0o ( OIollo0oLlLiI0IILOO00illIILLIoo0o ) , .O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ( O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ) , .OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ( OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ) , .OLli0lIO0lOO0OooILllIi00Lol00oili ( OLli0lIO0lOO0OooILllIi00Lol00oili ) , .Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ( Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ) , .OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ( OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ) , .OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ( OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ) , .OOIolooo0Oi00io00lIiiOiiLIliliOio ( OOIolooo0Oi00io00lIiiOiiLIliliOio ) , .OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ( OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ) , .O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ( O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ) , .OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ( OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ) , .OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ( OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ) , .Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ( Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ) , .O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ( O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ) , .OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ( OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ) , .OoI00LooIIlIIlIOOLIoloilI0OoIILLi ( OoI00LooIIlIIlIOOLIoloilI0OoIILLi ) , .OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ( OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ) , .O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ( O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ) , .OOIoOIilLi0looLILloOOollIIIo0llLo ( OOIoOIilLi0looLILloOOollIIIo0llLo ) , .OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ( OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ) , .OOllI0oo0L0io0l0IoloioOii0oIioOi0 ( OOllI0oo0L0io0l0IoloioOii0oIioOi0 ) , .OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ( OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ) , .Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ( Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ) , .O0oLiillllLOiLilOoI000iOLoiL0L0LO ( O0oLiillllLOiLilOoI000iOLoiL0L0LO ) , .OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ( OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ) , .Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ( Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ) , .OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ( OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ) , .OI0ioOlloiIio0oiOloi0lioiILoollLl ( OI0ioOlloiIio0oiOloi0lioiILoollLl ) , .OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ( OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ) , .OlIloooO00OIL0L0iIili0iOOoiLI0oiI ( OlIloooO00OIL0L0iIili0iOOoiLI0oiI ) , .OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ( OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ) , .OolIilIL0iooOLllOLloloOIlLIiOoLo0 ( OolIilIL0iooOLllOLloloOIlLIiOoLo0 ) , .OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ( OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ) , .OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ( OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ) , .O0lIOiilLOiIOollILlioiiOOiiLOO00i ( O0lIOiilLOiIOollILlioiiOOiiLOO00i ) , .O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ( O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ) , .OIiLIoliOIilIl0O00Li00oIO0OlIiooo ( OIiLIoliOIilIl0O00Li00oIO0OlIiooo ) , .OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ( OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ) , .O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ( O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ) , .Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ( Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ) , .Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ( Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ) , .OOoL0lOOloLLOLOILLLOolliIll0oOOoO ( OOoL0lOOloLLOLOILLLOolliIll0oOOoO ) , .OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ( OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ) , .OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ( OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ) , .O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ( O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ) , .OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ( OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ) , .O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ( O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ) , .O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ( O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ) , .OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ( OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ) , .OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ( OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ) , .Ol000OloII0LlIII00IIOIlOiioOo0Iii ( Ol000OloII0LlIII00IIOIlOiioOo0Iii ) , .OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ( OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ) , .OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ( OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ) , .OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ( OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ) , .OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ( OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ) , .OLLli0LLl0LlILOoi000iLoiiOOOLooLI ( OLLli0LLl0LlILOoi000iLoiiOOOLooLI ) , .OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ( OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ) , .OoooIiooOl0i0oliO0lio0IOo0iIILLLi ( OoooIiooOl0i0oliO0lio0IOo0iIILLLi ) , .OoOlILlliliiOI0OLLoOOl0000iIo0IIo ( OoOlILlliliiOI0OLLoOOl0000iIo0IIo ) , .OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ( OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ) , .O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ( O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ) , .OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ( OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ) , .OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ( OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ) , .OLolLol0lLIIlIillI000oIlilLLloOii ( OLolLol0lLIIlIillI000oIlilLLloOii ) , .OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ( OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ) , .OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ( OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ) , .OO0O0oOlliIoIOlooIO0lOLolIilLllIO ( OO0O0oOlliIoIOlooIO0lOLolIilLllIO ) , .O00I0iOoILll0oILl0ILloii0LIIOOiIO ( O00I0iOoILll0oILl0ILloii0LIIOOiIO ) , .OlolloloolOo0o0LLLIl00Li0iiLl00ol ( OlolloloolOo0o0LLLIl00Li0iiLl00ol ) , .OIIli0ilooIlOLI0lLO0Oi0IilILOolii ( OIIli0ilooIlOLI0lLO0Oi0IilILOolii ) , .OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ( OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ) , .OoOOLol000OllOLI0LO0LO0LoIliO0iiL ( OoOOLol000OllOLI0LO0LO0LoIliO0iiL ) , .OoIooi0LILolioIilliiol0I0iLoioIoi ( OoIooi0LILolioIilliiol0I0iLoioIoi ) , .OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ( OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ) , .OLlLoL0lO0oOIOolIIoiILIO0oOilooll ( OLlLoL0lO0oOIOolIIoiILIO0oOilooll ) , .O0iI0Lil0liLOLiILLOoilII0LII0iolO ( O0iI0Lil0liLOLiILLOoilII0LII0iolO ) , .OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ( OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ) , .OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ( OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ) , .O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ( O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ) , .OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ( OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ) , .OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ( OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ) , .OLLloO00IliLiLLlLloLloO0liOoIIOOI ( OLLloO00IliLiLLlLloLloO0liOoIIOOI ) , .OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ( OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ) , .OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ( OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ) , .OO00IIiOlOioiOLIiIloilLII0lLL0OOi ( OO00IIiOlOioiOLIiIloilLII0lLL0OOi ) , .OOLIlLlLIloIOoooilolooLloIi0OiiIi ( OOLIlLlLIloIOoooilolooLloIi0OiiIi ) , .OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ( OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ) , .OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ( OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ) , .OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ( OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ) , .OILolilliOIlLILOoioLii0iI0lII0oil ( OILolilliOIlLILOoioLii0iI0lII0oil ) , .OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ( OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ) , .OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ( OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ) , .O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ( O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ) , .OoLLliL00LLoooll00ooiLolOliOO0lLI ( OoLLliL00LLoooll00ooiLolOliOO0lLI ) , .OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ( OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ) , .O00loOoIIlII0OOo0lio00iOOOolLiIiO ( O00loOoIIlII0OOo0lio00iOOOolLiIiO ) , .OiiOIoolI0LioIo0IlL0lOllILIOOiIio ( OiiOIoolI0LioIo0IlL0lOllILIOOiIio ) , .OoIooolIllLIIolLII0IiLLiiOlOOIIOO ( OoIooolIllLIIolLII0IiLLiiOlOOIIOO ) , .OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ( OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ) , .OLL0i00LllLlio0oLOLooIL0ilLLllil0 ( OLL0i00LllLlio0oLOLooIL0ilLLllil0 ) , .OOiOiOIIoOii0oOLlI0OliIi0liioLLII ( OOiOiOIIoOii0oOLlI0OliIi0liioLLII ) , .OlOl0iOIioolOiill0OLOloOoLiIlllol ( OlOl0iOIioolOiill0OLOloOoLiIlllol ) , .OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ( OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ) , .OloILiOiLoIOOl0IoloOlI00Oollol0lL ( OloILiOiLoIOOl0IoloOlI00Oollol0lL ) , .OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ( OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ) , .OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ( OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ) , .OOIilioOiLLoOIL0iLoILiLLliiio0LOl ( OOIilioOiLLoOIL0iLoILiLLliiio0LOl ) , .O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ( O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ) , .Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ( Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ) , .O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ( O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ) , .O0li0llLIi0oIo0IilLLooLILolLIOOoo ( O0li0llLIi0oIo0IilLLooLILolLIOOoo ) , .OioIOIo0IllIo0OILLlli0LOOl00lioII ( OioIOIo0IllIo0OILLlli0LOOl00lioII ) , .OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ( OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ) , .OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ( OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ) , .Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ( Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ) , .OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ( OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ) , .OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ( OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ) , .O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ( O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ) , .OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ( OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ) , .OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ( OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ) , .O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ( O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ) , .OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ( OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ) , .OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ( OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ) , .OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ( OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ) , .OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ( OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ) , .Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ( Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ) , .O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ( O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ) , .OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ( OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ) , .O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ( O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ) , .O0il0OIIioo0IoL0OI0llOiLiLioill0i ( O0il0OIIioo0IoL0OI0llOiLiLioill0i ) , .O0lioOi00lO0IL00IoLLILolIlli00LiI ( O0lioOi00lO0IL00IoLLILolIlli00LiI ) , .OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ( OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ) , .OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ( OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ) , .OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ( OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ) , .OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ( OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ) , .OioOlIooLl0IL0LiioIlILIolO0o0ii0l ( OioOlIooLl0IL0LiioIlILIolO0o0ii0l ) , .OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ( OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ) , .OI0ILilL0olIiOoL0lOiiooolOOllIIIL ( OI0ILilL0olIiOoL0lOiiooolOOllIIIL ) , .O0000LloLiliiLOoIi0iLiLli0iloOOLI ( O0000LloLiliiLOoIi0iLiLli0iloOOLI ) , .OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ( OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ) , .OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ( OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ) , .OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ( OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ) , .OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ( OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ) , .OIO0IIi0OIooOiLOIII0lLolililiOIll ( OIO0IIi0OIooOiLOIII0lLolililiOIll ) , .OioilLoll0OiiOooiLiIOiL0LiilILII0 ( OioilLoll0OiiOooiLiIOiL0LiilILII0 ) , .OLoli0Li0i0oO0olOOilIliIio0LOoIIO ( OLoli0Li0i0oO0olOOilIliIio0LOoIIO ) , .OLLOoOIo0oiL0IOOO0lill0iloILllIOO ( OLLOoOIo0oiL0IOOO0lill0iloILllIOO ) , .OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ( OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ) , .OIILOOOOIOl00OoIollioiiliIilolLLl ( OIILOOOOIOl00OoIollioiiliIilolLLl ) , .OiooooLLoI0OLilIIil0ilooLo0OIloLl ( OiooooLLoI0OLilIIil0ilooLo0OIloLl ) , .O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ( O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ) , .OiLiiLILIoLilioiLolliOl0LI00LLil0 ( OiLiiLILIoLilioiLolliOl0LI00LLil0 ) , .Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ( Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ) , .Oloo0IIooolliliLOLoLoL0oI0LOliLlL ( Oloo0IIooolliliLOLoLoL0oI0LOliLlL ) , .OIiIIlooOiolooLoI0iLi0loLiloiLOll ( OIiIIlooOiolooLoI0iLi0loLiloiLOll ) , .OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ( OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ) , .OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ( OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ) , .OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ( OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ) , .OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ( OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ) , .Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ( Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ) , .OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ( OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ) , .Ol0OLoIiI0OloLIlillLOloLioIIL0III ( Ol0OLoIiI0OloLIlillLOloLioIIL0III ) , .OiILooool0OiolIOIIlO0LiOliIiIL0Ii ( OiILooool0OiolIOIIlO0LiOliIiIL0Ii ) , .OlLiiOLII0io0OLOOiIiiO0IIililoolo ( OlLiiOLII0io0OLOOiIiiO0IIililoolo ) , .OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ( OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ) , .OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ( OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ) , .OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ( OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ) , .OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ( OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ) , .OLlolloLliiLO0IlIlLo0lIiiloL00OOL ( OLlolloLliiLO0IlIlLo0lIiiloL00OOL ) , .OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ( OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ) , .O00oIiiOLOoilolOol0OIIOII00lllOIo ( O00oIiiOLOoilolOol0OIIOII00lllOIo ) , .OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ( OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ) , .OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ( OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ) , .Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ( Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ) , .OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ( OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ) , .OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ( OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ) , .OLi0ooOo0OlIllLOILllLL00lL00Liii0 ( OLi0ooOo0OlIllLOILllLL00lL00Liii0 ) , .OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ( OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ) , .Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ( Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ) , .OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ( OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ) , .Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ( Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ) , .Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ( Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ) , .OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ( OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ) , .OOOLilOolI0LILLIoloIiO00OiIiLiiIo ( OOOLilOolI0LILLIoloIiO00OiIiLiiIo ) , .OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ( OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ) , .OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ( OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ) , .OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ( OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ) , .OlLi0LOI0LoLioI0loilIlo00iliILIoi ( OlLi0LOI0LoLioI0loilIlo00iliILIoi ) , .OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ( OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ) , .OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ( OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ) , .OiOoiILoiIiIIoll0loilLl00Ll00O0iL ( OiOoiILoiIiIIoll0loilLl00Ll00O0iL ) , .OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ( OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ) , .OIlLiI0I0l0olLllLI0LliOOlllliLL0i ( OIlLiI0I0l0olLllLI0LliOOlllliLL0i ) , .OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ( OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ) , .OO0OOoLL0O0OOOllioILi0liilLLloiLO ( OO0OOoLL0O0OOOllioILi0liilLLloiLO ) , .OlLlliliOioioOIoiLOIOiOoiiioIOLOO ( OlLlliliOioioOIoiLOIOiOoiiioIOLOO ) , .OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ( OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ) , .OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ( OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ) , .OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ( OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ) , .OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ( OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ) , .OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ( OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ) , .OliliILl0LLiioool00L00LoLLILio0lO ( OliliILl0LLiioool00L00LoLLILio0lO ) , .OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ( OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ) , .OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ( OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ) , .OLioIOLOILilililoO0ililOi0oiIoo0o ( OLioIOLOILilililoO0ililOi0oiIoo0o ) , .OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ( OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ) , .Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ( Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ) , .Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ( Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ) , .OioIoIoo0iIIlOilLlIoILioo0I0lo00o ( OioIoIoo0iIIlOilLlIoILioo0I0lo00o ) , .O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ( O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ) , .OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ( OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ) , .OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ( OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ) , .OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ( OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ) , .O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ( O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ) , .OoLiLLooILIo0iol0OIoliLi0iiioiIlI ( OoLiLLooILIo0iol0OIoliLi0iiioiIlI ) , .OI0ool0i0ollOOoloL00L0LlLIO0LIliI ( OI0ool0i0ollOOoloL00L0LlLIO0LIliI ) , .Oo0loliLllliloIiliOi0lILloLI0ILlO ( Oo0loliLllliloIiliOi0lILloLI0ILlO ) , .Ooi0OL0i0IioliooLiI00OoiL00looOIL ( Ooi0OL0i0IioliooLiI00OoiL00looOIL ) , .OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ( OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ) , .OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ( OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ) , .OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ( OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ) , .OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ( OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ) , .OoOLolo0o0IOilOOLI0OoioLilIliI0lO ( OoOLolo0o0IOilOOLI0OoioLilIliI0lO ) , .O0o0OiliollLIi0IiLilIiOlLOOOLO00i ( O0o0OiliollLIi0IiLilIiOlLOOOLO00i ) , .OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ( OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ) , .OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ( OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ) , .OOIILlIiIOiOIi0o0li0lolol0LIoOliI ( OOIILlIiIOiOIi0o0li0lolol0LIoOliI ) , .OOIlIio0iILll00lliIIioiIiOLlLLi00 ( OOIlIio0iILll00lliIIioiIiOLlLLi00 ) , .OlIollIiLi0IlLiolloLOOL000Oo0l0II ( OlIollIiLi0IlLiolloLOOL000Oo0l0II ) , .OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ( OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ) , .OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ( OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ) , .OiiooiLLOL0iiO0oILoOlLoololiIIo0o ( OiiooiLLOL0iiO0oILoOlLoololiIIo0o ) , .OL0Lio0lIililolilllOL0Li0lIi0I0LI ( OL0Lio0lIililolilllOL0Li0lIi0I0LI ) , .O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ( O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ) , .OolL0oo00LOo0LOoLiILllLo0loOoIiii ( OolL0oo00LOo0LOoLiILllLo0loOoIiii ) , .OIOIOlilIolIlLOLlLlll0IiOIiILiOol ( OIOIOlilIolIlLOLlLlll0IiOIiILiOol ) , .OiloLLIlO00Il0oo0io0Iilliiil0OolO ( OiloLLIlO00Il0oo0io0Iilliiil0OolO ) , .O0oOL0illOloooo0ioIiOLOooLILllLl0 ( O0oOL0illOloooo0ioIiOLOooLILllLl0 ) , .Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ( Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ) , .OlOL0OLLooilLiOliIOIOOlIio00Oiili ( OlOL0OLLooilLiOliIOIOOlIio00Oiili ) , .OO0oolOlI0iloil0ooIolIioiol00I00I ( OO0oolOlI0iloil0ooIolIioiol00I00I ) , .O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ( O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ) , .OLI00Il0O0lI0OoLI0oIloiOIiiILIill ( OLI00Il0O0lI0OoLI0oIloiOIiiILIill ) , .OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ( OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ) , .OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ( OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ) , .O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ( O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ) , .OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ( OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ) , .OOoLol0oioL0looOlO0io0oIillil0iI0 ( OOoLol0oioL0looOlO0io0oIillil0iI0 ) , .OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ( OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ) , .OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ( OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ) , .O0oilLoOiOiLLi0Li0lLOIooIiliILlii ( O0oilLoOiOiLLi0Li0lLOIooIiliILlii ) , .O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ( O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ) , .OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ( OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ) , .OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ( OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ) , .OLiILioillIololIOILoOLlI0LILLliIL ( OLiILioillIololIOILoOLlI0LILLliIL ) , .OoOOillllIiloIOIILO0lL0LIl0iOlIII ( OoOOillllIiloIOIILO0lL0LIl0iOlIII ) , .OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ( OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ) , .OLIoIliI0LI0liL0i0IIIiLloL000l0lO ( OLIoIliI0LI0liL0i0IIIiLloL000l0lO ) , .Oo00OloiOIoLi00Oo0ooiololoOoooLLO ( Oo00OloiOIoLi00Oo0ooiololoOoooLLO ) , .Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ( Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ) , .Ollil0L0OlO0loio0OLiLILo0OioO0iOO ( Ollil0L0OlO0loio0OLiLILo0OioO0iOO ) , .OLio000LoL0lOol0oIiLlILLIlOLLOIlO ( OLio000LoL0lOol0oIiLlILLIlOLLOIlO ) , .OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ( OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ) , .OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ( OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ) , .OILIi00LOILOoLIiLloLiLIolliOoooIo ( OILIi00LOILOoLIiLloLiLIolliOoooIo ) , .OioilI0Oo0oOil0lIioiILIOLLLOLLioO ( OioilI0Oo0oOil0lIioiILIOLLLOLLioO ) , .OI0L0iIOilOi0LlILL0l0liiiil0lOIii ( OI0L0iIOilOi0LlILL0l0liiiil0lOIii ) , .OlIIioIIlILoli0oIiIl0l0IlOlloooll ( OlIIioIIlILoli0oIiIl0l0IlOlloooll ) , .O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ( O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ) , .OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ( OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ) , .OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ( OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ) , .Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ( Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ) , .OIOO0oiiIiiOILOOioiiO00OIl0lilllO ( OIOO0oiiIiiOILOOioiiO00OIl0lilllO ) , .OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ( OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ) , .OO0iLILOLioOioLOoLIOlOlo0oOIollll ( OO0iLILOLioOioLOoLIOlOlo0oOIollll ) , .OI00OlLIOIiOOiIliIooII00LLLllLLOO ( OI00OlLIOIiOOiIliIooII00LLLllLLOO ) , .OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ( OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ) , .O0L0O0ioooOOiLLlLLOLiioooILolII0o ( O0L0O0ioooOOiLLlLLOLiioooILolII0o ) , .OoiiooOo00OI0O0loiolLOLioIOiI0LoI ( OoiiooOo00OI0O0loiolLOLioIOiI0LoI ) , .OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ( OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ) , .O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ( O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ) , .OIi0liIIIoiOooLllLO0O0IoLLllIOlli ( OIi0liIIIoiOooLllLO0O0IoLLllIOlli ) , .OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ( OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ) , .OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ( OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ) , .OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ( OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ) , .OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ( OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ) , .OI0OLOILiOlOoolLIilooolollLLo0OOO ( OI0OLOILiOlOoolLIilooolollLLo0OOO ) , .O0Il0L0lLloiIiliL0000o0oIOLLILool ( O0Il0L0lLloiIiliL0000o0oIOLLILool ) , .OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ( OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ) , .Oo00IIIIoOIO0IL00llOoOioiollIOi00 ( Oo00IIIIoOIO0IL00llOoOioiollIOi00 ) , .OlIliOioiio0LLoLl00i0liioIOI00iIi ( OlIliOioiio0LLoLl00i0liioIOI00iIi ) , .OLOlLlooLIlL0IIiOilIiIooLloIioLOi ( OLOlLlooLIlL0IIiOilIiIooLloIioLOi ) , .OOlOiiLoIooll0L00oIIIoOIililiillo ( OOlOiiLoIooll0L00oIIIoOIililiillo ) , .O0i000LoOoll00lolOOOOIO0Oio0LIO0o ( O0i000LoOoll00lolOOOOIO0Oio0LIO0o ) , .OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ( OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ) , .Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ( Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ) , .OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ( OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ) , .O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ( O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ) , .O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ( O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ) , .O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ( O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ) , .OooOIi00Ii0liOollOoLioI0OiLiLiO0O ( OooOIi00Ii0liOollOoLioI0OiLiLiO0O ) , .OioolLOlII0IlolOIiLOliilL0oiiOoIo ( OioolLOlII0IlolOIiLOliilL0oiiOoIo ) , .OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ( OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ) , .OoII0il0iLlL00iIo0I0OoloiiilLOLIo ( OoII0il0iLlL00iIo0I0OoloiiilLOLIo ) , .OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ( OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ) , .Oi0Liloll0L00OiL0iLli0LO00iloIoLi ( Oi0Liloll0L00OiL0iLli0LO00iloIoLi ) , .OolIl0OOoiOlLioiloO0OolLOiIOolLLI ( OolIl0OOoiOlLioiloO0OolLOiIOolLLI ) , .OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ( OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ) , .OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ( OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ) , .OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ( OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ) , .Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ( Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ) , .OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ( OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ) , .OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ( OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ) , .O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ( O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ) , .OO0llOooLooLoi0l0oIOOoilOolIoLLOo ( OO0llOooLooLoi0l0oIOOoilOolIoLLOo ) , .OOIIlilOoOlIolLlILLioil0LL0oLlloo ( OOIIlilOoOlIolLlILLioil0LL0oLlloo ) , .OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ( OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ) , .OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ( OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ) , .OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ( OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ) , .OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ( OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ) , .Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ( Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ) , .OOoooLL0l0llOLI0o0oO00LIoLO00LILO ( OOoooLL0l0llOLI0o0oO00LIoLO00LILO ) , .OoilLIlliloO0LoOL00IILioiolLIloi0 ( OoilLIlliloO0LoOL00IILioiolLIloi0 ) , .OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ( OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ) , .O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ( O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ) , .OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ( OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ) , .Oll00iO0Ol0IOLloLLilo0OliIloIiLli ( Oll00iO0Ol0IOLloLLilo0OliIloIiLli ) , .OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ( OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ) , .OLllIIIO0oIlllOo00LILooILo0io0o00 ( OLllIIIO0oIlllOo00LILooILo0io0o00 ) , .OIO0IioIOoIOIll0LOIlOOILoILoiilli ( OIO0IioIOoIOIll0LOIlOOILoILoiilli ) , .Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ( Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ) , .OLl0oiiIOL0ol00LIoo0IoolIollol0ii ( OLl0oiiIOL0ol00LIoo0IoolIollol0ii ) , .OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ( OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ) , .OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ( OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ) , .OiILIII00lOolOiililIOiIIloo0OlLlo ( OiILIII00lOolOiililIOiIIloo0OlLlo ) , .OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ( OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ) , .OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ( OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ) , .OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ( OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ) , .OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ( OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ) , .OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ( OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ) , .O0lIi00lIl0iOlLilOloOIllllLLolooo ( O0lIi00lIl0iOlLilOloOIllllLLolooo ) , .OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ( OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ) , .O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ( O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ) , .OIl0iolIOLOlLOloIoLoIo0OooLi000lO ( OIl0iolIOLOlLOloIoLoIo0OooLi000lO ) , .Oiio0oo000ioIO0llioIoLILlIlIOOloL ( Oiio0oo000ioIO0llioIoLILlIlIOOloL ) , .OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ( OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ) , .OLoOLiILLLiIilOolo0Lil0iLLOOLILII ( OLoOLiILLLiIilOolo0Lil0iLLOOLILII ) , .O00liliooOOoiI0OlOOIIlO0o0IiOOolL ( O00liliooOOoiI0OlOOIIlO0o0IiOOolL ) , .OILLl0iillioLoOiiIiL0iliIOiO0oiio ( OILLl0iillioLoOiiIiL0iliIOiO0oiio ) , .OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ( OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ) , .O0I0LooLLiIO0illo0IliLLoioL0LlOLl ( O0I0LooLLiIO0illo0IliLLoioL0LlOLl ) , .OiioOooilOllI0oOoolilo0OLIlioo0II ( OiioOooilOllI0oOoolilo0OLIlioo0II ) , .OIolOIIiLIloloOL0iIIO0il0li00ilOo ( OIolOIIiLIloloOL0iIIO0il0li00ilOo ) , .OlOllIloiIIIIloliooOo0LoIil0o0oii ( OlOllIloiIIIIloliooOo0LoIil0o0oii ) , .OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ( OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ) , .OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ( OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ) , .OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ( OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ) , .OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ( OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ) , .OLILoOooIiil0oIIolILIlLIioL0i0Iio ( OLILoOooIiil0oIIolILIlLIioL0i0Iio ) , .OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ( OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ) , .OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ( OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ) , .OIooL0lILLIloiOOLiI0ilOIli0LOL000 ( OIooL0lILLIloiOOLiI0ilOIli0LOL000 ) , .O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ( O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ) , .OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ( OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ) , .O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ( O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ) , .OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ( OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ) , .OOiOiIiiilililLoLlIOoIoiILilLoooI ( OOiOiIiiilililLoLlIOoIoiILilLoooI ) , .OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ( OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ) , .OIiolOOI00iliL0LolLOOOLOliiIlLlII ( OIiolOOI00iliL0LolLOOOLOliiIlLlII ) , .O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ( O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ) , .O0OoiooiIOLOllil0OLoLOlllL000LII0 ( O0OoiooiIOLOllil0OLoLOlllL000LII0 ) , .Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ( Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ) , .OOl0i0OIIooLiI0IioL0LLILIloOlOllL ( OOl0i0OIIooLiI0IioL0LLILIloOlOllL ) , .OOOlLolILloIii0oollOil0lI0OOoOoo0 ( OOOlLolILloIii0oollOil0lI0OOoOoo0 ) , .O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ( O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ) , .O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ( O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ) , .OOI0llLoO0IOO000OilllLLLI0i0Iilil ( OOI0llLoO0IOO000OilllLLLI0i0Iilil ) , .OOIOl00lliliioILLoiioolL0OLLoLo0i ( OOIOl00lliliioILLoiioolL0OLLoLo0i ) , .OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ( OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ) , .OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ( OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ) , .OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ( OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ) , .Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ( Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ) , .OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ( OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ) , .OO0O00OIoioOIOLi0IlILI0OlilooOIOo ( OO0O00OIoioOIOLi0IlILI0OlilooOIOo ) , .OlLo00LioOiOOOoliolIoLI0olOOlLoOI ( OlLo00LioOiOOOoliolIoLI0olOOlLoOI ) , .OLOL0OioiLOLoli0LOL00OOiO0iiOooll ( OLOL0OioiLOLoli0LOL00OOiO0iiOooll ) , .OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ( OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ) , .O0oiOOLLiiillOliOOOllO0iO000OOoLI ( O0oiOOLLiiillOliOOOllO0iO000OOoLI ) , .OIliOOilOillIo00oiOOLIOiLolIIooOl ( OIliOOilOillIo00oiOOLIOiLolIIooOl ) , .OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ( OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ) , .OIlOIiiliIlIOIlilliilOl0iILIOOOLO ( OIlOIiiliIlIOIlilliilOl0iILIOOOLO ) , .OIoll0OLiliiLlIililii0oiII0Ol00lO ( OIoll0OLiliiLlIililii0oiII0Ol00lO ) , .Ol0LliIIIIiOOILo0ooioLolOOOololIo ( Ol0LliIIIIiOOILo0ooioLolOOOololIo ) , .OlollLLLoL0iiI0lool0OOOOIiOoolioL ( OlollLLLoL0iiI0lool0OOOOIiOoolioL ) , .O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ( O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ) , .OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ( OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ) , .OllloLIILloiiiOill0lOLooilli0Llii ( OllloLIILloiiiOill0lOLooilli0Llii ) , .OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ( OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ) , .OlLIiOlioIILOllO00lLiI0LiIlOloIiI ( OlLIiOlioIILOllO00lLiI0LiIlOloIiI ) , .OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ( OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ) , .OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ( OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ) , .OliiLi0oooOIo0L0lLoil0ooooi00I0ol ( OliiLi0oooOIo0L0lLoil0ooooi00I0ol ) , .O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ( O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ) , .OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ( OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ) , .OlIIloOL0iLIOLlOlLILlloiioloooILi ( OlIIloOL0iLIOLlOlLILlloiioloooILi ) , .OolOOLl0OlII0OiiloIloOO00IllliiLO ( OolOOLl0OlII0OiiloIloOO00IllliiLO ) , .O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ( O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ) , .OIliolloLooOi0OolOOi0ILOlIliLi0o0 ( OIliolloLooOi0OolOOi0ILOlIliLi0o0 ) , .Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ( Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ) , .OIILiOiLOO0IILI0llIOoooi0oLiiOioO ( OIILiOiLOO0IILI0llIOoooi0oLiiOioO ) , .OLOILIii00lILOLoLIIlOiioll0ilOLii ( OLOILIii00lILOLoLIIlOiioll0ilOLii ) , .O0IlliiI0l00iOLL0oLilIILo00lLIolo ( O0IlliiI0l00iOLL0oLilIILo00lLIolo ) , .OII0Iill0IOLO000li0iL0iLoiIoOoliL ( OII0Iill0IOLO000li0iL0iLoiIoOoliL ) , .OoIL0ll0llIOoI0IoIioiILILllLLOOOL ( OoIL0ll0llIOoI0IoIioiILILllLLOOOL ) , .OlIli0IolOiL0LoliLloo0olllliIiO0O ( OlIli0IolOiL0LoliLloo0olllliIiO0O ) , .OO00il0IO0lLoiilIo0ioiOiOOlLloioL ( OO00il0IO0lLoiilIo0ioiOiOOlLloioL ) , .OLoLOlol00olO0oo0LLlolI0OiLo0llLI ( OLoLOlol00olO0oo0LLlolI0OiLo0llLI ) , .OlIiO0llI0O0Li00OLIILiOLi00OiLioL ( OlIiO0llI0O0Li00OLIILiOLi00OiLioL ) , .OoL0LLOIlII0oLlloILillo0IOilOi0Il ( OoL0LLOIlII0oLlloILillo0IOilOi0Il ) , .OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ( OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ) , .OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ( OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ) , .OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ( OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ) , .O0o0OillO0LllooIiILLoilol0lii0liL ( O0o0OillO0LllooIiILLoilol0lii0liL ) , .OIO0L0iO0iLllOLILO0IoLliLolI00lLI ( OIO0L0iO0iLllOLILO0IoLliLolI00lLI ) , .OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ( OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ) , .OoOll0iOi0l0LiioLllOoliOoO00Lloil ( OoOll0iOi0l0LiioLllOoliOoO00Lloil ) , .OiIoioILioOLl0io00oiOiO0liliOlOoO ( OiIoioILioOLl0io00oiOiO0liliOlOoO ) , .OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ( OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ) , .OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ( OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ) , .OOI0I0II0oOOO0LiLoO0I00LloOllilIl ( OOI0I0II0oOOO0LiLoO0I00LloOllilIl ) , .OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ( OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ) , .OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ( OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ) , .OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ( OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ) , .OLolOilolLoloilIloOOiioIloiI0L0Lo ( OLolOilolLoloilIloOOiioIloiI0L0Lo ) , .O0lIlL0lLL00000ioioloooIoiiiioi00 ( O0lIlL0lLL00000ioioloooIoiiiioi00 ) , .Oioo00O0OIloLlOil00lLiI0oIOOOoIio ( Oioo00O0OIloLlOil00lLiI0oIOOOoIio ) , .O0oL00LOlilLooOoiil0oLL0iIillLlLL ( O0oL00LOlilLooOoiil0oLL0iIillLlLL ) , .OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ( OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ) , .OOILlooOIliLloiliIOi00LIlLIoli000 ( OOILlooOIliLloiliIOi00LIlLIoli000 ) , .OLOlILilLoI0liOiooL00OOlo0i0LiiiI ( OLOlILilLoI0liOiooL00OOlo0i0LiiiI ) , .O0oOLILIoIlLOIIollLOoL00o0O00OiOo ( O0oOLILIoIlLOIIollLOoL00o0O00OiOo ) , .O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ( O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ) , .OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ( OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ) , .O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ( O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ) , .O0OllOiIO00LliIOoLolo0loIiL0LiIlI ( O0OllOiIO00LliIOoLolo0loIiL0LiIlI ) , .OOOOLL0II0ioIiIIoLOolIOLIoLooIill ( OOOOLL0II0ioIiIIoLOolIOLIoLooIill ) , .OOIioIlLoOL00lOliIIllL00illo0L00o ( OOIioIlLoOL00lOliIIllL00illo0L00o ) , .OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ( OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ) , .Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ( Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ) , .O0oIiILIIO0LOOil00IlIoLiIilO00ooI ( O0oIiILIIO0LOOil00IlIoLiIilO00ooI ) , .OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ( OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ) , .OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ( OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ) , .OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ( OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ) , .Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ( Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ) , .OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ( OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ) , .OiIL00IOiOiiI00oiio0lLOlooIiLiOio ( OiIL00IOiOiiI00oiio0lLOlooIiLiOio ) , .OOIIilloi0OiOoo0iI0LI0LI00oILiLio ( OOIIilloi0OiOoo0iI0LI0LI00oILiLio ) , .Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ( Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ) , .OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ( OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ) , .O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ( O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ) , .Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ( Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ) , .Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ( Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ) , .OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ( OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ) , .OLiloooloollOoil0LlolLolOILlO00Ol ( OLiloooloollOoil0LlolLolOILlO00Ol ) , .O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ( O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ) , .OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ( OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ) , .OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ( OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ) , .OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ( OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ) , .OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ( OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ) , .O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ( O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ) , .OIOio00oLLL0o00LO00LLoI0LlL0OILlO ( OIOio00oLLL0o00LO00LLoI0LlL0OILlO ) , .OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ( OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ) , .O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ( O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ) , .OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ( OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ) , .OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ( OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ) , .O0illollo0oliIl0OolOoIlIILL0OIioO ( O0illollo0oliIl0OolOoIlIILL0OIioO ) , .O0Il00oIILloI0IL0LiOO0i0lIiIoolio ( O0Il00oIILloI0IL0LiOO0i0lIiIoolio ) , .OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ( OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ) , .OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ( OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ) , .OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ( OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ) , .OOilLILioilLIliOlOoilOOIolLLiLl0I ( OOilLILioilLIliOlOoilOOIolLLiLl0I ) , .OiOo0O0ooiioi00lloILL0oLLoILOiLiO ( OiOo0O0ooiioi00lloILL0oLLoILOiLiO ) , .OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ( OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ) , .OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ( OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ) , .OLololIl0LoiLooLIloiooLli0LOOLLli ( OLololIl0LoiLooLIloiooLli0LOOLLli ) , .OILllI0lillIoilOIoooOll0LII00I0l0 ( OILllI0lillIoilOIoooOll0LII00I0l0 ) , .OLiILL00lIlOliLloi0OOl00LlIl0Loli ( OLiILL00lIlOliLloi0OOl00LlIl0Loli ) , .OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ( OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ) , .OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ( OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ) , .OilIl00OOIloIli0LIIii00LIIlILiL0L ( OilIl00OOIloIli0LIIii00LIIlILiL0L ) , .OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ( OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ) , .OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ( OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ) , .OoOoIOoI0LILoIlIliLIioOooOOOIOoli ( OoOoIOoI0LILoIlIliLIioOooOOOIOoli ) , .OI00OLIIi0LioLLLLllooOiOl0iolOO0I ( OI00OLIIi0LioLLLLllooOiOl0iolOO0I ) , .OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ( OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ) , .OLIIl0o0liIOIooiOII0liO0oLllOI0oO ( OLIIl0o0liIOIooiOII0liO0oLllOI0oO ) , .OlOiOoL0i0i0L00OL00l00OOoL0OLILol ( OlOiOoL0i0i0L00OL00l00OOoL0OLILol ) , .OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ( OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ) , .OlLILiOolLl0ioiLiLlILiILLlIOllloI ( OlLILiOolLl0ioiLiLlILiILLlIOllloI ) , .OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ( OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ) , .OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ( OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ) , .OIllOIIOiOol000OoLIL0lLl0L00iIIIL ( OIllOIIOiOol000OoLIL0lLl0L00iIIIL ) , .OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ( OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ) , .OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ( OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ) , .OlLiolooLilLlLiil0l0iiO0IOILool00 ( OlLiolooLilLlLiil0l0iiO0IOILool00 ) , .OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ( OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ) , .OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ( OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ) , .OIoolOll00LlI00l0oIOLLIOI0I0LIILo ( OIoolOll00LlI00l0oIOLLIOI0I0LIILo ) , .OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ( OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ) , .OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ( OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ) , .OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ( OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ) , .OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ( OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ) , .Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ( Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ) , .OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ( OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ) , .OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ( OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ) , .OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ( OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ) , .O0lolLi0olIioIiIooOLLLlioIooLIill ( O0lolLi0olIioIiIooOLLLlioIooLIill ) , .OolLO0OOloooOIOiiOilL0IiILL0iol0I ( OolLO0OOloooOIOiiOilL0IiILL0iol0I ) , .OL0looio0Loioi0ill0olOo0o00ioOOII ( OL0looio0Loioi0ill0olOo0o00ioOOII ) , .Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ( Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ) , .Ol0LioliiiiOil0liLiOiolioOo0oioii ( Ol0LioliiiiOil0liLiOiolioOo0oioii ) , .Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ( Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ) , .OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ( OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ) , .OO0oIOllioLiLlLLlii0ilL0OlIliIilO ( OO0oIOllioLiLlLLlii0ilL0OlIliIilO ) , .OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ( OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ) , .OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ( OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ) , .OLOllOoI0IolOloolLolO0lIiolLiIILi ( OLOllOoI0IolOloolLolO0lIiolLiIILi ) , .OOILLooOOlllIILoIiIioLIOI0LOiLiLI ( OOILLooOOlllIILoIiIioLIOI0LOiLiLI ) , .O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ( O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ) , .OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ( OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ) , .Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ( Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ) , .OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ( OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ) , .O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ( O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ) , .OilO0OLOo0LllI00o0oOil00L0OloIOl0 (OilO0OLOo0LllI00o0oOil00L0OloIOl0 ) , .OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll (OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll ) , .OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l (OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l ) , .OILLiiO0o00OloIOOl0LlIOOlo00O0OOi (OILLiiO0o00OloIOOl0LlIOOlo00O0OOi ) , .OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil (OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil ) , .Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 (Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 ) , .OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl (OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl ) , .Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI (Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI ) , .OlolI00LoLoOILILoioLOL0lolLO0oiOo ( OlolI00LoLoOILILoioLOL0lolLO0oiOo ) , .OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL ( OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL ) , .O0000Lil0OoOOILlIlOlooioiIOloOioi ( O0000Lil0OoOOILlIlOlooioiIOloOioi ) , .O00lOOl0oILIoiioLOOI0OoioILioLiiL ( O00lOOl0oILIoiioLOOI0OoioILioLiiL ) , .O0iioiILo0ol0ollLilLl0lO0oI0ilOiL ( O0iioiILo0ol0ollLilLl0lO0oI0ilOiL ) );
 reg OllL0ooOlllIIOOi0iOOlIL0ol0I0IiOL;
 reg [255:0] Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL;
 reg [255:0] OiIOI0OLOLlliILOL0IoOLlLolil0OiIi;
 wire O0LOIOil0oI0OOOlOiILiLL0L0lLIOoIo;
 wire Oi00OiOiio0ILo00lL0lO0iLOOlIIOLLo;
 wire [255:0] OILoOilIOILLlOOLliI0oLlOoOIooolO0;
 wire [255:0] O0oOilLliiOiOi0O0I0llILlLoI0loLio = { OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 7: 0], OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 15: 8],OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 23: 16],OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 31: 24], OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 39: 32], OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 47: 40],OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 55: 48],OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 63: 56], OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 71: 64], OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 79: 72],OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 87: 80],OilO0OLOo0LllI00o0oOil00L0OloIOl0[ 95: 88], OilO0OLOo0LllI00o0oOil00L0OloIOl0[103: 96], OilO0OLOo0LllI00o0oOil00L0OloIOl0[111:104],OilO0OLOo0LllI00o0oOil00L0OloIOl0[119:112],OilO0OLOo0LllI00o0oOil00L0OloIOl0[127:120], OilO0OLOo0LllI00o0oOil00L0OloIOl0[135:128], OilO0OLOo0LllI00o0oOil00L0OloIOl0[143:136],OilO0OLOo0LllI00o0oOil00L0OloIOl0[151:144],OilO0OLOo0LllI00o0oOil00L0OloIOl0[159:152], OilO0OLOo0LllI00o0oOil00L0OloIOl0[167:160], OilO0OLOo0LllI00o0oOil00L0OloIOl0[175:168],OilO0OLOo0LllI00o0oOil00L0OloIOl0[183:176],OilO0OLOo0LllI00o0oOil00L0OloIOl0[191:184], OilO0OLOo0LllI00o0oOil00L0OloIOl0[199:192], OilO0OLOo0LllI00o0oOil00L0OloIOl0[207:200],OilO0OLOo0LllI00o0oOil00L0OloIOl0[215:208],OilO0OLOo0LllI00o0oOil00L0OloIOl0[223:216], OilO0OLOo0LllI00o0oOil00L0OloIOl0[231:224], OilO0OLOo0LllI00o0oOil00L0OloIOl0[239:232],OilO0OLOo0LllI00o0oOil00L0OloIOl0[247:240],OilO0OLOo0LllI00o0oOil00L0OloIOl0[255:248] };
 wire [255:0] OoOli0LiLl0LiO0olOI0IOoolliloIiO0 = { OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 7: 0], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 15: 8],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 23: 16],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 31: 24], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 39: 32], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 47: 40],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 55: 48],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 63: 56], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 71: 64], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 79: 72],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 87: 80],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[ 95: 88], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[103: 96], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[111:104],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[119:112],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[127:120], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[135:128], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[143:136],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[151:144],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[159:152], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[167:160], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[175:168],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[183:176],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[191:184], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[199:192], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[207:200],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[215:208],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[223:216], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[231:224], OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[239:232],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[247:240],OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll[255:248] };
 wire [255:0] O0ooLlOl0iLiIlOLlIIIIiol0IOL0iilo = { OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 7: 0], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 15: 8],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 23: 16],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 31: 24], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 39: 32], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 47: 40],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 55: 48],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 63: 56], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 71: 64], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 79: 72],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 87: 80],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[ 95: 88], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[103: 96], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[111:104],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[119:112],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[127:120], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[135:128], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[143:136],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[151:144],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[159:152], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[167:160], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[175:168],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[183:176],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[191:184], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[199:192], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[207:200],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[215:208],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[223:216], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[231:224], OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[239:232],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[247:240],OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil[255:248] };
 wire [255:0] OilIlI0IiI0LlLOiOLi00o0liOIiLLI0O = { Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 7: 0], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 15: 8],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 23: 16],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 31: 24], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 39: 32], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 47: 40],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 55: 48],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 63: 56], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 71: 64], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 79: 72],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 87: 80],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[ 95: 88], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[103: 96], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[111:104],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[119:112],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[127:120], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[135:128], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[143:136],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[151:144],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[159:152], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[167:160], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[175:168],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[183:176],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[191:184], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[199:192], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[207:200],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[215:208],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[223:216], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[231:224], Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[239:232],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[247:240],Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0[255:248] };
 wire [255:0] OiiLolOLLIii000ilOiIL0L0LILL0IILl = { OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 7: 0], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 15: 8],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 23: 16],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 31: 24], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 39: 32], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 47: 40],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 55: 48],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 63: 56], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 71: 64], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 79: 72],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 87: 80],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[ 95: 88], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[103: 96], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[111:104],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[119:112],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[127:120], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[135:128], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[143:136],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[151:144],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[159:152], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[167:160], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[175:168],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[183:176],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[191:184], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[199:192], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[207:200],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[215:208],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[223:216], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[231:224], OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[239:232],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[247:240],OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL[255:248] };
 wire [255:0] OiiIOlLl00loio0ioi00OlOLOoOllLLoI = { O0000Lil0OoOOILlIlOlooioiIOloOioi[ 7: 0], O0000Lil0OoOOILlIlOlooioiIOloOioi[ 15: 8],O0000Lil0OoOOILlIlOlooioiIOloOioi[ 23: 16],O0000Lil0OoOOILlIlOlooioiIOloOioi[ 31: 24], O0000Lil0OoOOILlIlOlooioiIOloOioi[ 39: 32], O0000Lil0OoOOILlIlOlooioiIOloOioi[ 47: 40],O0000Lil0OoOOILlIlOlooioiIOloOioi[ 55: 48],O0000Lil0OoOOILlIlOlooioiIOloOioi[ 63: 56], O0000Lil0OoOOILlIlOlooioiIOloOioi[ 71: 64], O0000Lil0OoOOILlIlOlooioiIOloOioi[ 79: 72],O0000Lil0OoOOILlIlOlooioiIOloOioi[ 87: 80],O0000Lil0OoOOILlIlOlooioiIOloOioi[ 95: 88], O0000Lil0OoOOILlIlOlooioiIOloOioi[103: 96], O0000Lil0OoOOILlIlOlooioiIOloOioi[111:104],O0000Lil0OoOOILlIlOlooioiIOloOioi[119:112],O0000Lil0OoOOILlIlOlooioiIOloOioi[127:120], O0000Lil0OoOOILlIlOlooioiIOloOioi[135:128], O0000Lil0OoOOILlIlOlooioiIOloOioi[143:136],O0000Lil0OoOOILlIlOlooioiIOloOioi[151:144],O0000Lil0OoOOILlIlOlooioiIOloOioi[159:152], O0000Lil0OoOOILlIlOlooioiIOloOioi[167:160], O0000Lil0OoOOILlIlOlooioiIOloOioi[175:168],O0000Lil0OoOOILlIlOlooioiIOloOioi[183:176],O0000Lil0OoOOILlIlOlooioiIOloOioi[191:184], O0000Lil0OoOOILlIlOlooioiIOloOioi[199:192], O0000Lil0OoOOILlIlOlooioiIOloOioi[207:200],O0000Lil0OoOOILlIlOlooioiIOloOioi[215:208],O0000Lil0OoOOILlIlOlooioiIOloOioi[223:216], O0000Lil0OoOOILlIlOlooioiIOloOioi[231:224], O0000Lil0OoOOILlIlOlooioiIOloOioi[239:232],O0000Lil0OoOOILlIlOlooioiIOloOioi[247:240],O0000Lil0OoOOILlIlOlooioiIOloOioi[255:248] };
 wire [31:0] O0oLlLIliIIOl0lI0iI0OiIlOIoiIliiO = { O00lOOl0oILIoiioLOOI0OoioILioLiiL[ 7: 0], O00lOOl0oILIoiioLOOI0OoioILioLiiL[ 15: 8],O00lOOl0oILIoiioLOOI0OoioILioLiiL[ 23: 16],O00lOOl0oILIoiioLOOI0OoioILioLiiL[ 31: 24] };
 reg [1:0] OILIIl0oOOoLooIIIi00I00L0ioOioo0L = 2'b0;
 always@ ( posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) OllL0ooOlllIIOOi0iOOlIL0ol0I0IiOL <= O0iioiILo0ol0ollLilLl0lO0oI0ilOiL;
 assign O0LOIOil0oI0OOOlOiILiLL0L0lLIOoIo = OllL0ooOlllIIOOi0iOOlIL0ol0I0IiOL ;
 always@ ( posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(O0iioiILo0ol0ollLilLl0lO0oI0ilOiL) OILIIl0oOOoLooIIIi00I00L0ioOioo0L <= OILIIl0oOOoLooIIIi00I00L0ioOioo0L + 1'b1;
 always@ ( posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(O0iioiILo0ol0ollLilLl0lO0oI0ilOiL && (OILIIl0oOOoLooIIIi00I00L0ioOioo0L == 2'b0) ) begin
 if(OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= O0oOilLliiOiOi0O0I0llILlLoI0loLio;
 else if(OILLiiO0o00OloIOOl0LlIOOlo00O0OOi) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= OoOli0LiLl0LiO0olOI0IOoolliloIiO0;
 else if(OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= O0ooLlOl0iLiIlOLlIIIIiol0IOL0iilo;
 else if(Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= OilIlI0IiI0LlLOiOLi00o0liOIiLLI0O;
 end
 else if(O0iioiILo0ol0ollLilLl0lO0oI0ilOiL && (OILIIl0oOOoLooIIIi00I00L0ioOioo0L == 2'b1)) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= OiiLolOLLIii000ilOiIL0L0LILL0IILl;
 else if(O0iioiILo0ol0ollLilLl0lO0oI0ilOiL && (OILIIl0oOOoLooIIIi00I00L0ioOioo0L == 2'd2)) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= OiiIOlLl00loio0ioi00OlOLOoOllLLoI;
 else if(O0iioiILo0ol0ollLilLl0lO0oI0ilOiL && (OILIIl0oOOoLooIIIi00I00L0ioOioo0L == 2'd3)) Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL <= O0oLlLIliIIOl0lI0iI0OiIlOIoiIliiO;
 always@ ( posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) OlLlOiIi0OoLiIlI0OO0loo0o0lOo0oIi <= 1'b0;
 else OlLlOiIi0OoLiIlI0OO0loo0o0lOo0oIi <= O0LOIOil0oI0OOOlOiILiLL0L0lLIOoIo;
 always@ ( posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) OL0O0lL0lIILiOLLil0LoIIIlILLO00ll <= Oll0oiolLoLloiILOoOLlOLLLlIIoOIIL ;
 assign OLlLLIloIliiIloOLloolLoIlLoi0iIoO = 1'd0 ;
 /* */ /* */ endmodule
 module OlLIO0oiil0ooIiOOioiLOI0oooilILoi ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI , OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 , OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol , OloliIooiiLI0IIlOiL0LLlioILLllL0L , O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO , OioILlIiO0000OoolooO00loIOIloLIoI , OLOl0000OLooLIIo0lIOIOI0lILioolOl , OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII , OoIolLlOIIoIoi00lloLlIoI0lo0iILol , OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI , OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo , OOIIloOlOILliIOILOIOiIlooIOOIL0oO , OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io , OiLOo0loOI00OL0Ooio0OIIlOLiooLOII , OlLilll0ilOLI0IIoO0li0l0OlO00oLIO , O0liLooiLliIoLOllliIlo0ILo0I0oOOl , O0i00oOl00OoIIOIil0LLOi0looIOIL00 , OlllLl0L0L0iO0lIloilOOo0iIIiOo00o , OOlOIlooi0LiIlLiilOL0LloiII0I0oLo , O0oLiillllLOiLilOoI000iOLoiL0L0LO , Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL , OoooIiooOl0i0oliO0lio0IOo0iIILLLi , OLlLoL0lO0oOIOolIIoiILIO0oOilooll , OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl , Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o , Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 , OLooLooiioOiOo00LLooO0OLoI0iLiLI0 , Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo , OLi0ooOo0OlIllLOILllLL00lL00Liii0 , OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I , OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o , OOIlIio0iILll00lliIIioiIiOLlLLi00 , OOiOLoILiiIiOLoOOOl0iOolLLloLLLil , OLio000LoL0lOol0oIiLlILLIlOLLOIlO , OoiiooOo00OI0O0loiolLOLioIOiI0LoI , Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl , OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I , OIO0IioIOoIOIll0LOIlOOILoILoiilli , OLoOLiILLLiIilOolo0Lil0iLLOOLILII , OOoLoi0LlLLLoIIllLLLIli0OI0LlliII , OiLl00LLioIio0iLiOiIOOOlLIlilOIOi , OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 , OlIli0IolOiL0LoliLloo0olllliIiO0O , OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 , Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 , OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO , OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 , OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo , O0lolLi0olIioIiIooOLLLlioIooLIill , OoolLolOioLILoOIII00LIOli00LIlloi , OOIolooo0Oi00io00lIiiOiiLIliliOio , OLLIiolLOOOliIoiIi0oLLiOllooIoiiI , OOoL0lOOloLLOLOILLLOolliIll0oOOoO , OoOlILlliliiOI0OLLoOOl0000iIo0IIo , O0iI0Lil0liLOLiILLOoilII0LII0iolO , O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 , O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI , O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 , OIO0IIi0OIooOiLOIII0lLolililiOIll , OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 , OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl , OO0OOoLL0O0OOOllioILi0liilLLloiLO , OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 , OlIollIiLi0IlLiolloLOOL000Oo0l0II , O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO , OOoIIOoIl0LIOllIO0L0oLoOIOoooiill , OiOIOlILOi0lIoOiIOIoOIllLILLiIliL , OO0LO0iliiL0Oi0OIIloILLOiO0LLloli , O00OiooIolIi0oIoIiiLlO0IiIO0ooLio , Oo0i0IlILOo0ooOiIlLOoiioll0LilllO , O00liliooOOoiI0OlOOIIlO0o0IiOOolL , O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI , Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO , OlLIiOlioIILOllO00lLiI0LiIlOloIiI , OO00il0IO0lLoiilIo0ioiOiOOlLloioL , OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl , O0oIiILIIO0LOOil00IlIoLiIilO00ooI , OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l , OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 , OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 , OolLO0OOloooOIOiiOilL0IiILL0iol0I , OOOooLlOLO0iOOOLi00oIiloILlooOLIO , OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI , Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi , OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO , OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO , OlL0ioloIOIoOLILilIIlIiLo0oIliOLI , OoLLliL00LLoooll00ooiLolOliOO0lLI , O0li0llLIi0oIo0IilLLooLILolLIOOoo , OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl , OioilLoll0OiiOooiLiIOiL0LiilILII0 , Ol0OLoIiI0OloLIlillLOloLioIIL0III , Oi0lll0000oiiLo0lOolIi0ooOiiI0lio , OlLlliliOioioOIoiLOIOiOoiiioIOLOO , OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 , OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO , OoIIiLoIL0llOo00oIi0oLi00oiill0Ll , OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili , O0IIL0iIliIIolLLiioLIILlIoI0o0IOI , O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO , OO0llOooLooLoi0l0oIOOoilOolIoLLOo , OLl0oiiIOL0ol00LIoo0IoolIollol0ii , OILLl0iillioLoOiiIiL0iliIOiO0oiio , OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 , OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 , OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I , OLoLOlol00olO0oo0LLlolI0OiLo0llLI , OLolOilolLoloilIloOOiioIloiI0L0Lo , OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi , OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o , OLololIl0LoiLooLIloiooLli0LOOLLli , OIllOIIOiOol000OoLIL0lLl0L00iIIIL , OL0looio0Loioi0ill0olOo0o00ioOOII , OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o , O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi , OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi , OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 , O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO , OLLIool0I0IooOOIoliL0Oo0iL0L0lOol , OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi , OioIOIo0IllIo0OILLlli0LOOl00lioII , O0l0lloOLloIiI0o0LIoi0LOllOIlO0io , OLoli0Li0i0oO0olOOilIliIio0LOoIIO , OiILooool0OiolIOIIlO0LiOliIiIL0Ii , OLIIoIiliIoiioIoLoI0LllolIIlO0LOi , OIlI0I0IooLOLIlLLLIlli0o0LLl0illI , O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 , OLLiIlIOlII00l00l0LoLLilL0l0OOOLo , OOoLol0oioL0looOlO0io0oIillil0iI0 , OILIi00LOILOoLIiLloLiLIolliOoooIo , OIi0liIIIoiOooLllLO0O0IoLLllIOlli , O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI , OOIIlilOoOlIolLlILLioil0LL0oLlloo , OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 , OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL , OOiOiIiiilililLoLlIOoIoiILilLoooI , OO0O00OIoioOIOLi0IlILI0OlilooOIOo , OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO , OlIiO0llI0O0Li00OLIILiOLi00OiLioL , O0lIlL0lLL00000ioioloooIoiiiioi00 , OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 , OioLlLLli0IiOllll0l0LiIoLiLLLOL0L , OILllI0lillIoilOIoooOll0LII00I0l0 , OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL , Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI , OioLioLloIiilLLoOlIoiLIO0IOoiLoll , OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo , OI0ioOlloiIio0oiOloi0lioiILoollLl , O0L0Ll0OOOO0O0oLloilIliooOLlILoIL , OiL0l0OlOOOLiOIliO0lII0OliliioOo0 , O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l , O00loOoIIlII0OOo0lio00iOOOolLiIiO , OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI , O0il0OIIioo0IoL0OI0llOiLiLioill0i , OLLOoOIo0oiL0IOOO0lill0iloILllIOO , OlLiiOLII0io0OLOOiIiiO0IIililoolo , Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO , OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 , OoLiLLooILIo0iol0OIoliLi0iiioiIlI , OiiooiLLOL0iiO0oILoOlLoololiIIo0o , OOlILLi0LIOoLiill0I0LOIOiOLoOO00I , OioilI0Oo0oOil0lIioiILIOLLLOLLioO , OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I , O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi , OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo , OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi , O0I0LooLLiIO0illo0IliLLoioL0LlOLl , OliI0i0iIOiOoiII0olii0OOO0LIOiLLi , OlLo00LioOiOOOoliolIoLI0olOOlLoOI , OliiLi0oooOIo0L0lLoil0ooooi00I0ol , OoL0LLOIlII0oLlloILillo0IOilOi0Il , Oioo00O0OIloLlOil00lLiI0oIOOOoIio , OIoOOO00OOolil0OIiIlllOOOo0Oil0oo , O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL , OLiILL00lIlOliLloi0OOl00LlIl0Loli , OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli , Ol0LioliiiiOil0liLiOiolioOo0oioii , Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi , OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi , OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO , OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL , OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI , OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 , OiiOIoolI0LioIo0IlL0lOllILIOOiIio , OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l , O0lioOi00lO0IL00IoLLILolIlli00LiI , OOiiIi0oILLIllilLLLOiIi0Ii0lii0II , OoiOoio0IOIoOio0olOLllllOIlLIoiL0 , Oi00i0oL0iIiLll0o0o0l0loi000ioOOL , OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo , OI0ool0i0ollOOoloL00L0LlLIO0LIliI , OL0Lio0lIililolilllOL0Li0lIi0I0LI , OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 , OI0L0iIOilOi0LlILL0l0liiiil0lOIii , OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL , OooOIi00Ii0liOollOoLioI0OiLiLiO0O , OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol , OiILIII00lOolOiililIOiIIloo0OlLlo , OiioOooilOllI0oOoolilo0OLIlioo0II , OIiolOOI00iliL0LolLOOOLOliiIlLlII , OLOL0OioiLOLoli0LOL00OOiO0iiOooll , O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO , OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo , O0oL00LOlilLooOoiil0oLL0iIillLlLL , Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl , OIOio00oLLL0o00LO00LLoI0LlL0OILlO , OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 , OlLiolooLilLlLiil0l0iiO0IOILool00 , Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i , OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 , Oo000ooL0O00L0illOlOLOO0oilOIi0Ll , OlIloooO00OIL0L0iIili0iOOoiLI0oiI , O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL , OLolLol0lLIIlIillI000oIlilLLloOii , OoIoIO0O0oOoilLlI000OIllIIoI0ioIl , OoIooolIllLIIolLII0IiLLiiOlOOIIOO , Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio , OI0i0lOolo0oOILo00ll0LIIOiOOlIoii , OIILOOOOIOl00OoIollioiiliIilolLLl , OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 , OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L , OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L , Oo0loliLllliloIiliOi0lILloLI0ILlO , O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io , O0oilLoOiOiLLi0Li0lLOIooIiliILlii , OlIIioIIlILoli0oIiIl0l0IlOlloooll , OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO , OioolLOlII0IlolOIiLOliilL0oiiOoIo , OLIoilIIoI0Ol0Oll0I0LloliiLlolIII , OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 , OIolOIIiLIloloOL0iIIO0il0li00ilOo , O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO , OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L , OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl , OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL , OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L , OIL0OiIiiiOLliIioloLo0lLILolLoLL0 , OILLLoLI0LiOLilloOiLOIlILI0Io0l0o , OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl , OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI , OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 , OIiO0OLioLiIOIIiLoiLooI00I0olI00O , O0Ol0i0loLlooOIiLoOlIilLolOlio0ll , OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I , O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi , OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo , OLLloO00IliLiLLlLloLloO0liOoIIOOI , OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi , OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI , OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L , OiooooLLoI0OLilIIil0ilooLo0OIloLl , OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO , OOOLilOolI0LILLIoloIiO00OiIiLiiIo , OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l , Ooi0OL0i0IioliooLiI00OoiL00looOIL , OolL0oo00LOo0LOoLiILllLo0loOoIiii , O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l , O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I , OllLlOiLLooiILOiiOOlLlL0LOII0LLOL , OilO0i0Lll00Iolo00lOOLiLiOiLO0lio , OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 , OLOl00iiILoiI00i0lOlLOi00IOLLlOIL , OlOllIloiIIIIloliooOo0LoIil0o0oii , O0OoiooiIOLOllil0OLoLOlllL000LII0 , O0oiOOLLiiillOliOOOllO0iO000OOoLI , OlIIloOL0iLIOLlOlLILlloiioloooILi , OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l , OOILlooOIliLloiliIOi00LIlLIoli000 , OiIL00IOiOiiI00oiio0lLOlooIiLiOio , O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo , OilIl00OOIloIli0LIIii00LIIlILiL0L , OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I , OO0oIOllioLiLlLLlii0ilL0OlIliIilO , OOOo0I0LlloiIl0i0il0OLiOlooOOolil , OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li , OolIilIL0iooOLllOLloloOIlLIiOoLo0 , OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO , OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 , OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl , OLL0i00LllLlio0oLOLooIL0ilLLllil0 , OLLLllOIlLOioiIIoOIOiLOILOioLlLLo , OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I , O0iooIILOi0llLIIoILoo0ilIIIlooLI0 , OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 , OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl , OliliILl0LLiioool00L00LoLLILio0lO , OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O , OIOIOlilIolIlLOLlLlll0IiOIiILiOol , OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo , OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 , OI0OLOILiOlOoolLIilooolollLLo0OOO , OoII0il0iLlL00iIo0I0OoloiiilLOLIo , Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l , OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl , OLIoLi0ioO0OLLl0LlIOillIoili0OIOI , Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i , OIliOOilOillIo00oiOOLIOiLolIIooOl , OolOOLl0OlII0OiiloIloOO00IllliiLO , O0o0OillO0LllooIiILLoilol0lii0liL , OLOlILilLoI0liOiooL00OOlo0i0LiiiI , OOIIilloi0OiOoo0iI0LI0LI00oILiLio , OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 , OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O , OIoolOll00LlI00l0oIOLLIOI0I0LIILo , OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 , OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o , OoI00LooIIlIIlIOOLIoloilI0OoIILLi , OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII , OL0OIiOoo0IllO0oloolIll0oOo0LlIIi , OO0O0oOlliIoIOlooIO0lOLolIilLllIO , OOIlLIiol0o00OlI0lLl0lILiIolL0iIi , OOiOiOIIoOii0oOLlI0OliIi0liioLLII , O0oiILoiiI0oOOoiillLOoiIilI0o0Ool , OI0O0lOIO0OOOOllIL00Ooi0I0llLlili , OiLiiLILIoLilioiLolliOl0LI00LLil0 , OLlolloLliiLO0IlIlLo0lIiiloL00OOL , OooLI0lioLIOiOOI00oLLOiLIOlO00ILi , OL0Oloi0OoLOiO00LLloIolIo0iiLLOII , OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo , OiloLLIlO00Il0oo0io0Iilliiil0OolO , OLI0iO0OLLO00l00LIlOLiiLlloILOLIl , OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I , O0Il0L0lLloiIiliL0000o0oIOLLILool , OiI0ILIIIiiLO0LOlOLliioLL0II0OooL , OOoooLL0l0llOLI0o0oO00LIoLO00LILO , OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl , OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 , OOl0i0OIIooLiI0IioL0LLILIloOlOllL , OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO , O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O , OIO0L0iO0iLllOLILO0IoLliLolI00lLI , O0oOLILIoIlLOIIollLOoL00o0O00OiOo , Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl , OoooO0olOolLIIOLIIl0L0ooLIOoOOioL , OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o , OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 , OLoOO0OOIooLoI0liLOLllIiIOIL0Olol , OLlOlii00IoIl00oIioIiIool0lLiOoLo , OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL , OL0LLioOOooILOL0LLLIilLl0oLLiIoiL , Ol000OloII0LlIII00IIOIlOiioOo0Iii , O00I0iOoILll0oILl0ILloii0LIIOOiIO , OO00IIiOlOioiOLIiIloilLII0lLL0OOi , OlOl0iOIioolOiill0OLOloOoLiIlllol , OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 , OioOlIooLl0IL0LiioIlILIolO0o0ii0l , Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 , OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO , OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol , OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII , OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 , O0oOL0illOloooo0ioIiOLOooLILllLl0 , OLiILioillIololIOILoOLlI0LILLliIL , Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 , OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 , Oi0Liloll0L00OiL0iLli0LO00iloIoLi , OoilLIlliloO0LoOL00IILioiolLIloi0 , OLIloIl0iIiooOIo0lLlO0L00LOIil0LO , OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO , OOOlLolILloIii0oollOil0lI0OOoOoo0 , OIlOIiiliIlIOIlilliilOl0iILIOOOLO , OIliolloLooOi0OolOOi0ILOlIliLi0o0 , OI00OOL0LLOOLLLiIooi0oL0iioOloL0O , O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L , OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 , O0illollo0oliIl0OolOoIlIILL0OIioO , OoOoIOoI0LILoIlIliLIioOooOOOIOoli , OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L , OLOllOoI0IolOloolLolO0lIiolLiIILi , OIollo0oLlLiI0IILOO00illIILLIoo0o , O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 , O0lIOiilLOiIOollILlioiiOOiiLOO00i , OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I , OlolloloolOo0o0LLLIl00Li0iiLl00ol , OOLIlLlLIloIOoooilolooLloIi0OiiIi , OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO , OlIoO0LIi0LOLoLLOoliioiIOolIl00OO , OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI , Oloo0IIooolliliLOLoLoL0oI0LOliLlL , O00oIiiOLOoilolOol0OIIOII00lllOIo , OlLi0LOI0LoLioI0loilIlo00iliILIoi , OLioIOLOILilililoO0ililOi0oiIoo0o , OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL , Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo , OoOOillllIiloIOIILO0lL0LIl0iOlIII , OIOO0oiiIiiOILOOioiiO00OIl0lilllO , Oo00IIIIoOIO0IL00llOoOioiollIOi00 , OolIl0OOoiOlLioiloO0OolLOiIOolLLI , OL00oOoLi0iLl00LILOOLOlooiiLOOoLo , O0lIi00lIl0iOlLilOloOIllllLLolooo , OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL , O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 , OIoll0OLiliiLlIililii0oiII0Ol00lO , Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi , OoOll0iOi0l0LiioLllOoliOoO00Lloil , OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 , O00o0iOOoOiLI0iiIOoIiIliLoIliIIll , O0Il00oIILloI0IL0LiOO0i0lIiIoolio , OI00OLIIi0LioLLLLllooOiOl0iolOO0I , OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO , OOILLooOOlllIILoIiIioLIOI0LOiLiLI , O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL , OOIoOIilLi0looLILloOOollIIIo0llLo , O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL , OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll , OIIli0ilooIlOLI0lLO0Oi0IilILOolii , OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO , OloILiOiLoIOOl0IoloOlI00Oollol0lL , O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L , OI0ILilL0olIiOoL0lOiiooolOOllIIIL , OIiIIlooOiolooLoI0iLi0loLiloiLOll , OO0ilOiiOiIooOlIiO0l00iOliILoOIIi , OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO , OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL , OoOLolo0o0IOilOOLI0OoioLilIliI0lO , OlOL0OLLooilLiOliIOIOOlIio00Oiili , OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi , OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO , OlIliOioiio0LLoLl00i0liioIOI00iIi , OOiiILOoLlI00LoOil0OiOoIlloIiOi0o , O0ioLLo0liLOOiOL0OoLiOool0lLI00oi , OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o , OLILoOooIiil0oIIolILIlLIioL0i0Iio , O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O , Ol0LliIIIIiOOILo0ooioLolOOOololIo , OIILiOiLOO0IILI0llIOoooi0oLiiOioO , OiIoioILioOLl0io00oiOiO0liliOlOoO , O0OOOLLL0oOLoillIiOLIiIoI00LioiLl , Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo , OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO , OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO , OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO , O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi , OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi , OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL , OIiLIoliOIilIl0O00Li00oIO0OlIiooo , OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I , OlOlIILOLLIll0lo0lO0IOliliOOiL0oI , OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO , OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI , OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl , O0000LloLiliiLOoIi0iLiLli0iloOOLI , OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl , OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI , OI00ilIioiLo0ioiiIi0O0IolOiOi00IO , Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll , O0o0OiliollLIi0IiLilIiOlLOOOLO00i , OO0oolOlI0iloil0ooIolIioiol00I00I , OLIoIliI0LI0liL0i0IIIiLloL000l0lO , OO0iLILOLioOioLOoLIOlOlo0oOIollll , OLOlLlooLIlL0IIiOilIiIooLloIioLOi , OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 , OoIlL0lI0iL0iiIoLii0lLLio00lIIOol , O0O0L0iLLIlOILiOLoIiLiliiIllIi0li , OOLIlOoI0oOlII0oIllLi0l00iOioLIOi , OOI0llLoO0IOO000OilllLLLI0i0Iilil , OlollLLLoL0iiI0lool0OOOOIiOoolioL , OLOILIii00lILOLoLIIlOiioll0ilOLii , OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol , O0OllOiIO00LliIOoLolo0loIiL0LiIlI , Ooo00lolOl0OIoLOIlIliL0oLooIolLiL , OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol , OLIIl0o0liIOIooiOII0liO0oLllOI0oO , Olo0llLLi0L0IiLooLi0IooLOol0iIiIO , OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O , OLli0lIO0lOO0OooILllIi00Lol00oili , OOllI0oo0L0io0l0IoloioOii0oIioOi0 , OIIli0o0iiLOoOlilIoLIooOIooIL0ilI , OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio , OoOOLol000OllOLI0LO0LO0LoIliO0iiL , OoLOolIOLlOIIlIiOioiIIOL0lioliOIi , OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI , OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo , OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil , OI0IOio0lIIOiLllLLLIoIoiIoiOLillO , Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI , OiOoiILoiIiIIoll0loilLl00Ll00O0iL , Oo0IoILIliiOo0oooOLOiIo00i0L00Iio , OOooiloOoOIIiOiiLlLlLlIOIOIlolIol , O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI , Oo00OloiOIoLi00Oo0ooiololoOoooLLO , OI00OlLIOIiOOiIliIooII00LLLllLLOO , OOlOiiLoIooll0L00oIIIoOIililiillo , OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 , Oll00iO0Ol0IOLloLLilo0OliIloIiLli , OIl0iolIOLOlLOloIoLoIo0OooLi000lO , OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI , OOIOl00lliliioILLoiioolL0OLLoLo0i , O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 , O0IlliiI0l00iOLL0oLilIILo00lLIolo , OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl , OOOOLL0II0ioIiIIoLOolIOLIoLooIill , OLLI0ilo0LiioOLloOLloiioiIoOiLl0O , OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO , OlOiOoL0i0i0L00OL00l00OOoL0OLILol , OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO , Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l , Ooii00l0ooOoIliILL0lLLLLLoILlIIoO , OILl0LOii0lOi0LlLIIoIL0LLOoli0oll , O0Io0oIliooLo0i0i0lL0IlILOloiiIlI , OLLli0LLl0LlILOoi000iLoiiOOOLooLI , OoIooi0LILolioIilliiol0I0iLoioIoi , OILolilliOIlLILOoioLii0iI0lII0oil , OOIilioOiLLoOIL0iLoILiLLliiio0LOl , OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l , OllioLi0iLLoIOlILoIL0oOO0OiIliOOi , OlOoOLLlO0LOilOiiOoiOi0o0lollolLl , OILoioOioIOL0lIOLoIlIOlolLiOLlIoo , OoI0i0iiiL0ililIOLiL0IioLIL0IooOo , OioIoIoo0iIIlOilLlIoILioo0I0lo00o , OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 , OLI00Il0O0lI0OoLI0oIloiOIiiILIill , Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL , OioOiiiOlioLLOllo0IiIOiOOli0oi0LI , O0i000LoOoll00lolOOOOIO0Oio0LIO0o , Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO , OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl , Oiio0oo000ioIO0llioIoLILlIlIOOloL , OIooL0lILLIloiOOLiI0ilOIli0LOL000 , OILlOiiL00II0oiOlOoOI0lI00I0oIIIi , OLoOiiL00iolo0LOliOll0I0ILIOL0iLI , OII0Iill0IOLO000li0iL0iLoiIoOoliL , OOI0I0II0oOOO0LiLoO0I00LloOllilIl , OOIioIlLoOL00lOliIIllL00illo0L00o , OLiloooloollOoil0LlolLolOILlO00Ol , OOilLILioilLIliOlOoilOOIolLLiLl0I , OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 , OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI , OIiLOlOll0ol0OOLIo0oOiIilII0Io00L , OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI , Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO , Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi , OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI , OloIioIl0OOlolI0LIiioiLoL0OL0iI0i , OLIIoil00iiOOl0oloiiooOiI0IlL00Ol , O0L0oo0LI0OiII0l00oioIIiiilLLIOIl , OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl , OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo , OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI , OOoo0oiIolLIlol0oll00LiolIOOIlLL0 , OIlLiI0I0l0olLllLI0LliOOlllliLL0i , O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o , OOIILlIiIOiOIi0o0li0lolol0LIoOliI , OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL , Ollil0L0OlO0loio0OLiLILo0OioO0iOO , O0L0O0ioooOOiLLlLLOLiioooILolII0o , OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl , OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 , OLllIIIO0oIlllOo00LILooILo0io0o00 , OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI , O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO , OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 , OllloLIILloiiiOill0lOLooilli0Llii , OoIL0ll0llIOoI0IoIioiILILllLLOOOL , OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll , OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL , O0oLLI0O0IlOllolLIioIIOll0iiiIlLL , OiOo0O0ooiioi00lloILL0oLLoILOiLiO , OlLILiOolLl0ioiLiLlILiILLlIOllloI , OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O , O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi , OilO0OLOo0LllI00o0oOil00L0OloIOl0 , OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll , OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l , OILLiiO0o00OloIOOl0LlIOOlo00O0OOi , OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil , Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 , OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl , Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI , OlolI00LoLoOILILoioLOL0lolLO0oiOo , OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL , O0000Lil0OoOOILlIlOlooioiIOloOioi , O00lOOl0oILIoiioLOOI0OoioILioLiiL , O0iioiILo0ol0ollLilLl0lO0oI0ilOiL );
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 input [ 23: 0] OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI ;
 input [ 7: 0] OilIL0OIOillLolooIl0LLIo0lIL0Ooo0 ;
 input [ 31: 0] OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol ;
 input [ 7: 0] OloliIooiiLI0IIlOiL0LLlioILLllL0L ;
 input [ 31: 0] O0oLOOoILlLLoOIi0L0IiiillIOoL0oiO ;
 input [175: 0] OioILlIiO0000OoolooO00loIOIloLIoI ;
 input [ 71: 0] OLOl0000OLooLIIo0lIOIOI0lILioolOl ;
 input [ 31: 0] OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII ;
 input [ 63: 0] OoIolLlOIIoIoi00lloLlIoI0lo0iILol ;
 input [ 31: 0] OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI ;
 input [ 63: 0] OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo ;
 input [ 63: 0] OOIIloOlOILliIOILOIOiIlooIOOIL0oO ;
 input [ 63: 0] OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io ;
 input [ 31: 0] OiLOo0loOI00OL0Ooio0OIIlOLiooLOII ;
 input [ 63: 0] OlLilll0ilOLI0IIoO0li0l0OlO00oLIO ;
 input [ 31: 0] O0liLooiLliIoLOllliIlo0ILo0I0oOOl ;
 input O0i00oOl00OoIIOIil0LLOi0looIOIL00 ;
 input [ 23: 0] OlllLl0L0L0iO0lIloilOOo0iIIiOo00o ;
 input [ 23: 0] OOlOIlooi0LiIlLiilOL0LloiII0I0oLo ;
 input [ 23: 0] O0oLiillllLOiLilOoI000iOLoiL0L0LO ;
 input [ 23: 0] Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL ;
 input [ 23: 0] OoooIiooOl0i0oliO0lio0IOo0iIILLLi ;
 input [ 23: 0] OLlLoL0lO0oOIOolIIoiILIO0oOilooll ;
 input [ 23: 0] OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl ;
 input [ 23: 0] Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o ;
 input [ 23: 0] Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0 ;
 input [ 23: 0] OLooLooiioOiOo00LLooO0OLoI0iLiLI0 ;
 input [ 23: 0] Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo ;
 input [ 23: 0] OLi0ooOo0OlIllLOILllLL00lL00Liii0 ;
 input [ 23: 0] OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I ;
 input [ 23: 0] OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o ;
 input [ 23: 0] OOIlIio0iILll00lliIIioiIiOLlLLi00 ;
 input [ 23: 0] OOiOLoILiiIiOLoOOOl0iOolLLloLLLil ;
 input [ 23: 0] OLio000LoL0lOol0oIiLlILLIlOLLOIlO ;
 input [ 23: 0] OoiiooOo00OI0O0loiolLOLioIOiI0LoI ;
 input [ 23: 0] Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl ;
 input [ 23: 0] OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I ;
 input [ 23: 0] OIO0IioIOoIOIll0LOIlOOILoILoiilli ;
 input [ 23: 0] OLoOLiILLLiIilOolo0Lil0iLLOOLILII ;
 input [ 23: 0] OOoLoi0LlLLLoIIllLLLIli0OI0LlliII ;
 input [ 23: 0] OiLl00LLioIio0iLiOiIOOOlLIlilOIOi ;
 input [ 23: 0] OiOO0LOLIOO0LOlloIOIillolO0iIo0I0 ;
 input [ 23: 0] OlIli0IolOiL0LoliLloo0olllliIiO0O ;
 input [ 23: 0] OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0 ;
 input [ 23: 0] Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0 ;
 input [ 23: 0] OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO ;
 input [ 23: 0] OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0 ;
 input [ 23: 0] OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo ;
 input [ 23: 0] O0lolLi0olIioIiIooOLLLlioIooLIill ;
 input [ 7: 0] OoolLolOioLILoOIII00LIOli00LIlloi ;
 input [ 7: 0] OOIolooo0Oi00io00lIiiOiiLIliliOio ;
 input [ 7: 0] OLLIiolLOOOliIoiIi0oLLiOllooIoiiI ;
 input [ 7: 0] OOoL0lOOloLLOLOILLLOolliIll0oOOoO ;
 input [ 7: 0] OoOlILlliliiOI0OLLoOOl0000iIo0IIo ;
 input [ 7: 0] O0iI0Lil0liLOLiILLOoilII0LII0iolO ;
 input [ 7: 0] O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0 ;
 input [ 7: 0] O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI ;
 input [ 7: 0] O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0 ;
 input [ 7: 0] OIO0IIi0OIooOiLOIII0lLolililiOIll ;
 input [ 7: 0] OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0 ;
 input [ 7: 0] OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl ;
 input [ 7: 0] OO0OOoLL0O0OOOllioILi0liilLLloiLO ;
 input [ 7: 0] OlL0IOLIoOoilLoIIolLIILoLLI0i0I00 ;
 input [ 7: 0] OlIollIiLi0IlLiolloLOOL000Oo0l0II ;
 input [ 7: 0] O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO ;
 input [ 7: 0] OOoIIOoIl0LIOllIO0L0oLoOIOoooiill ;
 input [ 7: 0] OiOIOlILOi0lIoOiIOIoOIllLILLiIliL ;
 input [ 7: 0] OO0LO0iliiL0Oi0OIIloILLOiO0LLloli ;
 input [ 7: 0] O00OiooIolIi0oIoIiiLlO0IiIO0ooLio ;
 input [ 7: 0] Oo0i0IlILOo0ooOiIlLOoiioll0LilllO ;
 input [ 7: 0] O00liliooOOoiI0OlOOIIlO0o0IiOOolL ;
 input [ 7: 0] O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI ;
 input [ 7: 0] Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO ;
 input [ 7: 0] OlLIiOlioIILOllO00lLiI0LiIlOloIiI ;
 input [ 7: 0] OO00il0IO0lLoiilIo0ioiOiOOlLloioL ;
 input [ 7: 0] OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl ;
 input [ 7: 0] O0oIiILIIO0LOOil00IlIoLiIilO00ooI ;
 input [ 7: 0] OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l ;
 input [ 7: 0] OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0 ;
 input [ 7: 0] OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00 ;
 input [ 7: 0] OolLO0OOloooOIOiiOilL0IiILL0iol0I ;
 input [ 31: 0] OOOooLlOLO0iOOOLi00oIiloILlooOLIO ;
 input [ 31: 0] OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI ;
 input [ 31: 0] Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi ;
 input [ 31: 0] OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO ;
 input [ 31: 0] OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO ;
 input [ 31: 0] OlL0ioloIOIoOLILilIIlIiLo0oIliOLI ;
 input [ 31: 0] OoLLliL00LLoooll00ooiLolOliOO0lLI ;
 input [ 31: 0] O0li0llLIi0oIo0IilLLooLILolLIOOoo ;
 input [ 31: 0] OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl ;
 input [ 31: 0] OioilLoll0OiiOooiLiIOiL0LiilILII0 ;
 input [ 31: 0] Ol0OLoIiI0OloLIlillLOloLioIIL0III ;
 input [ 31: 0] Oi0lll0000oiiLo0lOolIi0ooOiiI0lio ;
 input [ 31: 0] OlLlliliOioioOIoiLOIOiOoiiioIOLOO ;
 input [ 31: 0] OLoolO0oO0io0IiiiOIIIllllLOO0O0O0 ;
 input [ 31: 0] OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO ;
 input [ 31: 0] OoIIiLoIL0llOo00oIi0oLi00oiill0Ll ;
 input [ 31: 0] OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili ;
 input [ 31: 0] O0IIL0iIliIIolLLiioLIILlIoI0o0IOI ;
 input [ 31: 0] O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO ;
 input [ 31: 0] OO0llOooLooLoi0l0oIOOoilOolIoLLOo ;
 input [ 31: 0] OLl0oiiIOL0ol00LIoo0IoolIollol0ii ;
 input [ 31: 0] OILLl0iillioLoOiiIiL0iliIOiO0oiio ;
 input [ 31: 0] OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0 ;
 input [ 31: 0] OOoILooiOiiiIll0oOLLIIoO0oLolIIo0 ;
 input [ 31: 0] OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I ;
 input [ 31: 0] OLoLOlol00olO0oo0LLlolI0OiLo0llLI ;
 input [ 31: 0] OLolOilolLoloilIloOOiioIloiI0L0Lo ;
 input [ 31: 0] OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi ;
 input [ 31: 0] OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o ;
 input [ 31: 0] OLololIl0LoiLooLIloiooLli0LOOLLli ;
 input [ 31: 0] OIllOIIOiOol000OoLIL0lLl0L00iIIIL ;
 input [ 31: 0] OL0looio0Loioi0ill0olOo0o00ioOOII ;
 input [ 7: 0] OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o ;
 input [ 7: 0] O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi ;
 input [ 7: 0] OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi ;
 input [ 7: 0] OOllIIoLLLooiiOoLiIi0loOO0ilO00O0 ;
 input [ 7: 0] O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO ;
 input [ 7: 0] OLLIool0I0IooOOIoliL0Oo0iL0L0lOol ;
 input [ 7: 0] OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi ;
 input [ 7: 0] OioIOIo0IllIo0OILLlli0LOOl00lioII ;
 input [ 7: 0] O0l0lloOLloIiI0o0LIoi0LOllOIlO0io ;
 input [ 7: 0] OLoli0Li0i0oO0olOOilIliIio0LOoIIO ;
 input [ 7: 0] OiILooool0OiolIOIIlO0LiOliIiIL0Ii ;
 input [ 7: 0] OLIIoIiliIoiioIoLoI0LllolIIlO0LOi ;
 input [ 7: 0] OIlI0I0IooLOLIlLLLIlli0o0LLl0illI ;
 input [ 7: 0] O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0 ;
 input [ 7: 0] OLLiIlIOlII00l00l0LoLLilL0l0OOOLo ;
 input [ 7: 0] OOoLol0oioL0looOlO0io0oIillil0iI0 ;
 input [ 7: 0] OILIi00LOILOoLIiLloLiLIolliOoooIo ;
 input [ 7: 0] OIi0liIIIoiOooLllLO0O0IoLLllIOlli ;
 input [ 7: 0] O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI ;
 input [ 7: 0] OOIIlilOoOlIolLlILLioil0LL0oLlloo ;
 input [ 7: 0] OLiiOLILl0LIlL00OlL0Oili00IiIlIl0 ;
 input [ 7: 0] OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL ;
 input [ 7: 0] OOiOiIiiilililLoLlIOoIoiILilLoooI ;
 input [ 7: 0] OO0O00OIoioOIOLi0IlILI0OlilooOIOo ;
 input [ 7: 0] OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO ;
 input [ 7: 0] OlIiO0llI0O0Li00OLIILiOLi00OiLioL ;
 input [ 7: 0] O0lIlL0lLL00000ioioloooIoiiiioi00 ;
 input [ 7: 0] OIioLLolLoll0iO0LoLo0ILlii0ilO0o0 ;
 input [ 7: 0] OioLlLLli0IiOllll0l0LiIoLiLLLOL0L ;
 input [ 7: 0] OILllI0lillIoilOIoooOll0LII00I0l0 ;
 input [ 7: 0] OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL ;
 input [ 7: 0] Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI ;
 input [ 31: 0] OioLioLloIiilLLoOlIoiLIO0IOoiLoll ;
 input [ 31: 0] OOOLLiI0l0IIL0OI0L0LOiIOLi0L0LOIo ;
 input [ 31: 0] OI0ioOlloiIio0oiOloi0lioiILoollLl ;
 input [ 31: 0] O0L0Ll0OOOO0O0oLloilIliooOLlILoIL ;
 input [ 31: 0] OiL0l0OlOOOLiOIliO0lII0OliliioOo0 ;
 input [ 31: 0] O00oO0I0lLoiOOlOI0liloLOIL0ioIi0l ;
 input [ 31: 0] O00loOoIIlII0OOo0lio00iOOOolLiIiO ;
 input [ 31: 0] OlLoiiiIiiOilOLIIOlIlOLiOiiolILoI ;
 input [ 31: 0] O0il0OIIioo0IoL0OI0llOiLiLioill0i ;
 input [ 31: 0] OLLOoOIo0oiL0IOOO0lill0iloILllIOO ;
 input [ 31: 0] OlLiiOLII0io0OLOOiIiiO0IIililoolo ;
 input [ 31: 0] Ool0ilo0l0IIOII0IIiLOoOoLiOiOoOiO ;
 input [ 31: 0] OLi0OOiLI0oioOOLo0oOI0OiioIiLO0l0 ;
 input [ 31: 0] OoLiLLooILIo0iol0OIoliLi0iiioiIlI ;
 input [ 31: 0] OiiooiLLOL0iiO0oILoOlLoololiIIo0o ;
 input [ 31: 0] OOlILLi0LIOoLiill0I0LOIOiOLoOO00I ;
 input [ 31: 0] OioilI0Oo0oOil0lIioiILIOLLLOLLioO ;
 input [ 31: 0] OLoLlL0OOlIllIiIiOOL0OloOlI00iL0I ;
 input [ 31: 0] O0OL00iLlLOLOii0oLoiiOLlOIoiLoLIi ;
 input [ 31: 0] OIOIO0io0oiOlLlI00oIlOIILLLoIo0lo ;
 input [ 31: 0] OoiOOioLiiIOoL0Iol00IolIlIOi0ioLi ;
 input [ 31: 0] O0I0LooLLiIO0illo0IliLLoioL0LlOLl ;
 input [ 31: 0] OliI0i0iIOiOoiII0olii0OOO0LIOiLLi ;
 input [ 31: 0] OlLo00LioOiOOOoliolIoLI0olOOlLoOI ;
 input [ 31: 0] OliiLi0oooOIo0L0lLoil0ooooi00I0ol ;
 input [ 31: 0] OoL0LLOIlII0oLlloILillo0IOilOi0Il ;
 input [ 31: 0] Oioo00O0OIloLlOil00lLiI0oIOOOoIio ;
 input [ 31: 0] OIoOOO00OOolil0OIiIlllOOOo0Oil0oo ;
 input [ 31: 0] O0ii0ILOo0lIO0LIoLlLiILIOOLo0LLIL ;
 input [ 31: 0] OLiILL00lIlOliLloi0OOl00LlIl0Loli ;
 input [ 31: 0] OloIIiloO0Oo0oOlIoLI0iioO0ILOiLli ;
 input [ 31: 0] Ol0LioliiiiOil0liLiOiolioOo0oioii ;
 input [175: 0] Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi ;
 input [175: 0] OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi ;
 input [175: 0] OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO ;
 input [175: 0] OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL ;
 input [175: 0] OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI ;
 input [175: 0] OoIlLi0I0llOlo0lool0LO0O0LlLOILi0 ;
 input [175: 0] OiiOIoolI0LioIo0IlL0lOllILIOOiIio ;
 input [175: 0] OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l ;
 input [175: 0] O0lioOi00lO0IL00IoLLILolIlli00LiI ;
 input [175: 0] OOiiIi0oILLIllilLLLOiIi0Ii0lii0II ;
 input [175: 0] OoiOoio0IOIoOio0olOLllllOIlLIoiL0 ;
 input [175: 0] Oi00i0oL0iIiLll0o0o0l0loi000ioOOL ;
 input [175: 0] OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo ;
 input [175: 0] OI0ool0i0ollOOoloL00L0LlLIO0LIliI ;
 input [175: 0] OL0Lio0lIililolilllOL0Li0lIi0I0LI ;
 input [175: 0] OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0 ;
 input [175: 0] OI0L0iIOilOi0LlILL0l0liiiil0lOIii ;
 input [175: 0] OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL ;
 input [175: 0] OooOIi00Ii0liOollOoLioI0OiLiLiO0O ;
 input [175: 0] OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol ;
 input [175: 0] OiILIII00lOolOiililIOiIIloo0OlLlo ;
 input [175: 0] OiioOooilOllI0oOoolilo0OLIlioo0II ;
 input [175: 0] OIiolOOI00iliL0LolLOOOLOliiIlLlII ;
 input [175: 0] OLOL0OioiLOLoli0LOL00OOiO0iiOooll ;
 input [175: 0] O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO ;
 input [175: 0] OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo ;
 input [175: 0] O0oL00LOlilLooOoiil0oLL0iIillLlLL ;
 input [175: 0] Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl ;
 input [175: 0] OIOio00oLLL0o00LO00LLoI0LlL0OILlO ;
 input [175: 0] OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00 ;
 input [175: 0] OlLiolooLilLlLiil0l0iiO0IOILool00 ;
 input [175: 0] Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i ;
 input [ 71: 0] OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0 ;
 input [ 71: 0] Oo000ooL0O00L0illOlOLOO0oilOIi0Ll ;
 input [ 71: 0] OlIloooO00OIL0L0iIili0iOOoiLI0oiI ;
 input [ 71: 0] O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL ;
 input [ 71: 0] OLolLol0lLIIlIillI000oIlilLLloOii ;
 input [ 71: 0] OoIoIO0O0oOoilLlI000OIllIIoI0ioIl ;
 input [ 71: 0] OoIooolIllLIIolLII0IiLLiiOlOOIIOO ;
 input [ 71: 0] Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio ;
 input [ 71: 0] OI0i0lOolo0oOILo00ll0LIIOiOOlIoii ;
 input [ 71: 0] OIILOOOOIOl00OoIollioiiliIilolLLl ;
 input [ 71: 0] OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0 ;
 input [ 71: 0] OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L ;
 input [ 71: 0] OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L ;
 input [ 71: 0] Oo0loliLllliloIiliOi0lILloLI0ILlO ;
 input [ 71: 0] O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io ;
 input [ 71: 0] O0oilLoOiOiLLi0Li0lLOIooIiliILlii ;
 input [ 71: 0] OlIIioIIlILoli0oIiIl0l0IlOlloooll ;
 input [ 71: 0] OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO ;
 input [ 71: 0] OioolLOlII0IlolOIiLOliilL0oiiOoIo ;
 input [ 71: 0] OLIoilIIoI0Ol0Oll0I0LloliiLlolIII ;
 input [ 71: 0] OL0IOILllOOO0OIOL0000LoO0llOo0Lo0 ;
 input [ 71: 0] OIolOIIiLIloloOL0iIIO0il0li00ilOo ;
 input [ 71: 0] O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO ;
 input [ 71: 0] OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L ;
 input [ 71: 0] OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl ;
 input [ 71: 0] OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL ;
 input [ 71: 0] OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L ;
 input [ 71: 0] OIL0OiIiiiOLliIioloLo0lLILolLoLL0 ;
 input [ 71: 0] OILLLoLI0LiOLilloOiLOIlILI0Io0l0o ;
 input [ 71: 0] OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl ;
 input [ 71: 0] OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI ;
 input [ 71: 0] OI0oL0loOli0oOIo0oi0lLlolOOiooIo0 ;
 input [ 31: 0] OIiO0OLioLiIOIIiLoiLooI00I0olI00O ;
 input [ 31: 0] O0Ol0i0loLlooOIiLoOlIilLolOlio0ll ;
 input [ 31: 0] OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I ;
 input [ 31: 0] O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi ;
 input [ 31: 0] OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo ;
 input [ 31: 0] OLLloO00IliLiLLlLloLloO0liOoIIOOI ;
 input [ 31: 0] OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi ;
 input [ 31: 0] OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI ;
 input [ 31: 0] OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L ;
 input [ 31: 0] OiooooLLoI0OLilIIil0ilooLo0OIloLl ;
 input [ 31: 0] OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO ;
 input [ 31: 0] OOOLilOolI0LILLIoloIiO00OiIiLiiIo ;
 input [ 31: 0] OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l ;
 input [ 31: 0] Ooi0OL0i0IioliooLiI00OoiL00looOIL ;
 input [ 31: 0] OolL0oo00LOo0LOoLiILllLo0loOoIiii ;
 input [ 31: 0] O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l ;
 input [ 31: 0] O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I ;
 input [ 31: 0] OllLlOiLLooiILOiiOOlLlL0LOII0LLOL ;
 input [ 31: 0] OilO0i0Lll00Iolo00lOOLiLiOiLO0lio ;
 input [ 31: 0] OILi0IiLoLOllLioi0oiOlIILl0oiOoi0 ;
 input [ 31: 0] OLOl00iiILoiI00i0lOlLOi00IOLLlOIL ;
 input [ 31: 0] OlOllIloiIIIIloliooOo0LoIil0o0oii ;
 input [ 31: 0] O0OoiooiIOLOllil0OLoLOlllL000LII0 ;
 input [ 31: 0] O0oiOOLLiiillOliOOOllO0iO000OOoLI ;
 input [ 31: 0] OlIIloOL0iLIOLlOlLILlloiioloooILi ;
 input [ 31: 0] OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l ;
 input [ 31: 0] OOILlooOIliLloiliIOi00LIlLIoli000 ;
 input [ 31: 0] OiIL00IOiOiiI00oiio0lLOlooIiLiOio ;
 input [ 31: 0] O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo ;
 input [ 31: 0] OilIl00OOIloIli0LIIii00LIIlILiL0L ;
 input [ 31: 0] OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I ;
 input [ 31: 0] OO0oIOllioLiLlLLlii0ilL0OlIliIilO ;
 input [ 63: 0] OOOo0I0LlloiIl0i0il0OLiOlooOOolil ;
 input [ 63: 0] OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li ;
 input [ 63: 0] OolIilIL0iooOLllOLloloOIlLIiOoLo0 ;
 input [ 63: 0] OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO ;
 input [ 63: 0] OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00 ;
 input [ 63: 0] OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl ;
 input [ 63: 0] OLL0i00LllLlio0oLOLooIL0ilLLllil0 ;
 input [ 63: 0] OLLLllOIlLOioiIIoOIOiLOILOioLlLLo ;
 input [ 63: 0] OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I ;
 input [ 63: 0] O0iooIILOi0llLIIoILoo0ilIIIlooLI0 ;
 input [ 63: 0] OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0 ;
 input [ 63: 0] OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl ;
 input [ 63: 0] OliliILl0LLiioool00L00LoLLILio0lO ;
 input [ 63: 0] OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O ;
 input [ 63: 0] OIOIOlilIolIlLOLlLlll0IiOIiILiOol ;
 input [ 63: 0] OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo ;
 input [ 63: 0] OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0 ;
 input [ 63: 0] OI0OLOILiOlOoolLIilooolollLLo0OOO ;
 input [ 63: 0] OoII0il0iLlL00iIo0I0OoloiiilLOLIo ;
 input [ 63: 0] Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l ;
 input [ 63: 0] OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl ;
 input [ 63: 0] OLIoLi0ioO0OLLl0LlIOillIoili0OIOI ;
 input [ 63: 0] Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i ;
 input [ 63: 0] OIliOOilOillIo00oiOOLIOiLolIIooOl ;
 input [ 63: 0] OolOOLl0OlII0OiiloIloOO00IllliiLO ;
 input [ 63: 0] O0o0OillO0LllooIiILLoilol0lii0liL ;
 input [ 63: 0] OLOlILilLoI0liOiooL00OOlo0i0LiiiI ;
 input [ 63: 0] OOIIilloi0OiOoo0iI0LI0LI00oILiLio ;
 input [ 63: 0] OI00OlliiO0LlIIiOoIL0oooi0LloLLo0 ;
 input [ 63: 0] OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O ;
 input [ 63: 0] OIoolOll00LlI00l0oIOLLIOI0I0LIILo ;
 input [ 63: 0] OlO0LlOLl00IIOIOiilooOLo0liLiIOl0 ;
 input [ 31: 0] OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o ;
 input [ 31: 0] OoI00LooIIlIIlIOOLIoloilI0OoIILLi ;
 input [ 31: 0] OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII ;
 input [ 31: 0] OL0OIiOoo0IllO0oloolIll0oOo0LlIIi ;
 input [ 31: 0] OO0O0oOlliIoIOlooIO0lOLolIilLllIO ;
 input [ 31: 0] OOIlLIiol0o00OlI0lLl0lILiIolL0iIi ;
 input [ 31: 0] OOiOiOIIoOii0oOLlI0OliIi0liioLLII ;
 input [ 31: 0] O0oiILoiiI0oOOoiillLOoiIilI0o0Ool ;
 input [ 31: 0] OI0O0lOIO0OOOOllIL00Ooi0I0llLlili ;
 input [ 31: 0] OiLiiLILIoLilioiLolliOl0LI00LLil0 ;
 input [ 31: 0] OLlolloLliiLO0IlIlLo0lIiiloL00OOL ;
 input [ 31: 0] OooLI0lioLIOiOOI00oLLOiLIOlO00ILi ;
 input [ 31: 0] OL0Oloi0OoLOiO00LLloIolIo0iiLLOII ;
 input [ 31: 0] OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo ;
 input [ 31: 0] OiloLLIlO00Il0oo0io0Iilliiil0OolO ;
 input [ 31: 0] OLI0iO0OLLO00l00LIlOLiiLlloILOLIl ;
 input [ 31: 0] OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I ;
 input [ 31: 0] O0Il0L0lLloiIiliL0000o0oIOLLILool ;
 input [ 31: 0] OiI0ILIIIiiLO0LOlOLliioLL0II0OooL ;
 input [ 31: 0] OOoooLL0l0llOLI0o0oO00LIoLO00LILO ;
 input [ 31: 0] OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl ;
 input [ 31: 0] OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0 ;
 input [ 31: 0] OOl0i0OIIooLiI0IioL0LLILIloOlOllL ;
 input [ 31: 0] OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO ;
 input [ 31: 0] O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O ;
 input [ 31: 0] OIO0L0iO0iLllOLILO0IoLliLolI00lLI ;
 input [ 31: 0] O0oOLILIoIlLOIIollLOoL00o0O00OiOo ;
 input [ 31: 0] Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl ;
 input [ 31: 0] OoooO0olOolLIIOLIIl0L0ooLIOoOOioL ;
 input [ 31: 0] OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o ;
 input [ 31: 0] OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0 ;
 input [ 31: 0] OLoOO0OOIooLoI0liLOLllIiIOIL0Olol ;
 input [ 63: 0] OLlOlii00IoIl00oIioIiIool0lLiOoLo ;
 input [ 63: 0] OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL ;
 input [ 63: 0] OL0LLioOOooILOL0LLLIilLl0oLLiIoiL ;
 input [ 63: 0] Ol000OloII0LlIII00IIOIlOiioOo0Iii ;
 input [ 63: 0] O00I0iOoILll0oILl0ILloii0LIIOOiIO ;
 input [ 63: 0] OO00IIiOlOioiOLIiIloilLII0lLL0OOi ;
 input [ 63: 0] OlOl0iOIioolOiill0OLOloOoLiIlllol ;
 input [ 63: 0] OOooOoIiooIliiO0LoLiOlOoIlOOo00I0 ;
 input [ 63: 0] OioOlIooLl0IL0LiioIlILIolO0o0ii0l ;
 input [ 63: 0] Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0 ;
 input [ 63: 0] OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO ;
 input [ 63: 0] OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol ;
 input [ 63: 0] OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII ;
 input [ 63: 0] OoLO0LoiiIL0lilol0oloO0loiLLiIIl0 ;
 input [ 63: 0] O0oOL0illOloooo0ioIiOLOooLILllLl0 ;
 input [ 63: 0] OLiILioillIololIOILoOLlI0LILLliIL ;
 input [ 63: 0] Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0 ;
 input [ 63: 0] OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0 ;
 input [ 63: 0] Oi0Liloll0L00OiL0iLli0LO00iloIoLi ;
 input [ 63: 0] OoilLIlliloO0LoOL00IILioiolLIloi0 ;
 input [ 63: 0] OLIloIl0iIiooOIo0lLlO0L00LOIil0LO ;
 input [ 63: 0] OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO ;
 input [ 63: 0] OOOlLolILloIii0oollOil0lI0OOoOoo0 ;
 input [ 63: 0] OIlOIiiliIlIOIlilliilOl0iILIOOOLO ;
 input [ 63: 0] OIliolloLooOi0OolOOi0ILOlIliLi0o0 ;
 input [ 63: 0] OI00OOL0LLOOLLLiIooi0oL0iioOloL0O ;
 input [ 63: 0] O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L ;
 input [ 63: 0] OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0 ;
 input [ 63: 0] O0illollo0oliIl0OolOoIlIILL0OIioO ;
 input [ 63: 0] OoOoIOoI0LILoIlIliLIioOooOOOIOoli ;
 input [ 63: 0] OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L ;
 input [ 63: 0] OLOllOoI0IolOloolLolO0lIiolLiIILi ;
 input [ 63: 0] OIollo0oLlLiI0IILOO00illIILLIoo0o ;
 input [ 63: 0] O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0 ;
 input [ 63: 0] O0lIOiilLOiIOollILlioiiOOiiLOO00i ;
 input [ 63: 0] OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I ;
 input [ 63: 0] OlolloloolOo0o0LLLIl00Li0iiLl00ol ;
 input [ 63: 0] OOLIlLlLIloIOoooilolooLloIi0OiiIi ;
 input [ 63: 0] OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO ;
 input [ 63: 0] OlIoO0LIi0LOLoLLOoliioiIOolIl00OO ;
 input [ 63: 0] OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI ;
 input [ 63: 0] Oloo0IIooolliliLOLoLoL0oI0LOliLlL ;
 input [ 63: 0] O00oIiiOLOoilolOol0OIIOII00lllOIo ;
 input [ 63: 0] OlLi0LOI0LoLioI0loilIlo00iliILIoi ;
 input [ 63: 0] OLioIOLOILilililoO0ililOi0oiIoo0o ;
 input [ 63: 0] OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL ;
 input [ 63: 0] Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo ;
 input [ 63: 0] OoOOillllIiloIOIILO0lL0LIl0iOlIII ;
 input [ 63: 0] OIOO0oiiIiiOILOOioiiO00OIl0lilllO ;
 input [ 63: 0] Oo00IIIIoOIO0IL00llOoOioiollIOi00 ;
 input [ 63: 0] OolIl0OOoiOlLioiloO0OolLOiIOolLLI ;
 input [ 63: 0] OL00oOoLi0iLl00LILOOLOlooiiLOOoLo ;
 input [ 63: 0] O0lIi00lIl0iOlLilOloOIllllLLolooo ;
 input [ 63: 0] OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL ;
 input [ 63: 0] O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0 ;
 input [ 63: 0] OIoll0OLiliiLlIililii0oiII0Ol00lO ;
 input [ 63: 0] Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi ;
 input [ 63: 0] OoOll0iOi0l0LiioLllOoliOoO00Lloil ;
 input [ 63: 0] OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0 ;
 input [ 63: 0] O00o0iOOoOiLI0iiIOoIiIliLoIliIIll ;
 input [ 63: 0] O0Il00oIILloI0IL0LiOO0i0lIiIoolio ;
 input [ 63: 0] OI00OLIIi0LioLLLLllooOiOl0iolOO0I ;
 input [ 63: 0] OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO ;
 input [ 63: 0] OOILLooOOlllIILoIiIioLIOI0LOiLiLI ;
 input [ 63: 0] O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL ;
 input [ 63: 0] OOIoOIilLi0looLILloOOollIIIo0llLo ;
 input [ 63: 0] O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL ;
 input [ 63: 0] OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll ;
 input [ 63: 0] OIIli0ilooIlOLI0lLO0Oi0IilILOolii ;
 input [ 63: 0] OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO ;
 input [ 63: 0] OloILiOiLoIOOl0IoloOlI00Oollol0lL ;
 input [ 63: 0] O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L ;
 input [ 63: 0] OI0ILilL0olIiOoL0lOiiooolOOllIIIL ;
 input [ 63: 0] OIiIIlooOiolooLoI0iLi0loLiloiLOll ;
 input [ 63: 0] OO0ilOiiOiIooOlIiO0l00iOliILoOIIi ;
 input [ 63: 0] OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO ;
 input [ 63: 0] OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL ;
 input [ 63: 0] OoOLolo0o0IOilOOLI0OoioLilIliI0lO ;
 input [ 63: 0] OlOL0OLLooilLiOliIOIOOlIio00Oiili ;
 input [ 63: 0] OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi ;
 input [ 63: 0] OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO ;
 input [ 63: 0] OlIliOioiio0LLoLl00i0liioIOI00iIi ;
 input [ 63: 0] OOiiILOoLlI00LoOil0OiOoIlloIiOi0o ;
 input [ 63: 0] O0ioLLo0liLOOiOL0OoLiOool0lLI00oi ;
 input [ 63: 0] OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o ;
 input [ 63: 0] OLILoOooIiil0oIIolILIlLIioL0i0Iio ;
 input [ 63: 0] O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O ;
 input [ 63: 0] Ol0LliIIIIiOOILo0ooioLolOOOololIo ;
 input [ 63: 0] OIILiOiLOO0IILI0llIOoooi0oLiiOioO ;
 input [ 63: 0] OiIoioILioOLl0io00oiOiO0liliOlOoO ;
 input [ 63: 0] O0OOOLLL0oOLoillIiOLIiIoI00LioiLl ;
 input [ 63: 0] Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo ;
 input [ 63: 0] OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO ;
 input [ 63: 0] OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO ;
 input [ 63: 0] OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO ;
 input [ 63: 0] O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi ;
 input [ 31: 0] OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi ;
 input [ 31: 0] OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL ;
 input [ 31: 0] OIiLIoliOIilIl0O00Li00oIO0OlIiooo ;
 input [ 31: 0] OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I ;
 input [ 31: 0] OlOlIILOLLIll0lo0lO0IOliliOOiL0oI ;
 input [ 31: 0] OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO ;
 input [ 31: 0] OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI ;
 input [ 31: 0] OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl ;
 input [ 31: 0] O0000LloLiliiLOoIi0iLiLli0iloOOLI ;
 input [ 31: 0] OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl ;
 input [ 31: 0] OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI ;
 input [ 31: 0] OI00ilIioiLo0ioiiIi0O0IolOiOi00IO ;
 input [ 31: 0] Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll ;
 input [ 31: 0] O0o0OiliollLIi0IiLilIiOlLOOOLO00i ;
 input [ 31: 0] OO0oolOlI0iloil0ooIolIioiol00I00I ;
 input [ 31: 0] OLIoIliI0LI0liL0i0IIIiLloL000l0lO ;
 input [ 31: 0] OO0iLILOLioOioLOoLIOlOlo0oOIollll ;
 input [ 31: 0] OLOlLlooLIlL0IIiOilIiIooLloIioLOi ;
 input [ 31: 0] OOl0oiloLLLIo0Li0ioloOiioLl0I00O0 ;
 input [ 31: 0] OoIlL0lI0iL0iiIoLii0lLLio00lIIOol ;
 input [ 31: 0] O0O0L0iLLIlOILiOLoIiLiliiIllIi0li ;
 input [ 31: 0] OOLIlOoI0oOlII0oIllLi0l00iOioLIOi ;
 input [ 31: 0] OOI0llLoO0IOO000OilllLLLI0i0Iilil ;
 input [ 31: 0] OlollLLLoL0iiI0lool0OOOOIiOoolioL ;
 input [ 31: 0] OLOILIii00lILOLoLIIlOiioll0ilOLii ;
 input [ 31: 0] OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol ;
 input [ 31: 0] O0OllOiIO00LliIOoLolo0loIiL0LiIlI ;
 input [ 31: 0] Ooo00lolOl0OIoLOIlIliL0oLooIolLiL ;
 input [ 31: 0] OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol ;
 input [ 31: 0] OLIIl0o0liIOIooiOII0liO0oLllOI0oO ;
 input [ 31: 0] Olo0llLLi0L0IiLooLi0IooLOol0iIiIO ;
 input [ 31: 0] OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O ;
 input [ 63: 0] OLli0lIO0lOO0OooILllIi00Lol00oili ;
 input [ 63: 0] OOllI0oo0L0io0l0IoloioOii0oIioOi0 ;
 input [ 63: 0] OIIli0o0iiLOoOlilIoLIooOIooIL0ilI ;
 input [ 63: 0] OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio ;
 input [ 63: 0] OoOOLol000OllOLI0LO0LO0LoIliO0iiL ;
 input [ 63: 0] OoLOolIOLlOIIlIiOioiIIOL0lioliOIi ;
 input [ 63: 0] OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI ;
 input [ 63: 0] OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo ;
 input [ 63: 0] OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil ;
 input [ 63: 0] OI0IOio0lIIOiLllLLLIoIoiIoiOLillO ;
 input [ 63: 0] Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI ;
 input [ 63: 0] OiOoiILoiIiIIoll0loilLl00Ll00O0iL ;
 input [ 63: 0] Oo0IoILIliiOo0oooOLOiIo00i0L00Iio ;
 input [ 63: 0] OOooiloOoOIIiOiiLlLlLlIOIOIlolIol ;
 input [ 63: 0] O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI ;
 input [ 63: 0] Oo00OloiOIoLi00Oo0ooiololoOoooLLO ;
 input [ 63: 0] OI00OlLIOIiOOiIliIooII00LLLllLLOO ;
 input [ 63: 0] OOlOiiLoIooll0L00oIIIoOIililiillo ;
 input [ 63: 0] OlIOlLIlLOIlLio00OIiLloIooIOo0ol0 ;
 input [ 63: 0] Oll00iO0Ol0IOLloLLilo0OliIloIiLli ;
 input [ 63: 0] OIl0iolIOLOlLOloIoLoIo0OooLi000lO ;
 input [ 63: 0] OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI ;
 input [ 63: 0] OOIOl00lliliioILLoiioolL0OLLoLo0i ;
 input [ 63: 0] O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0 ;
 input [ 63: 0] O0IlliiI0l00iOLL0oLilIILo00lLIolo ;
 input [ 63: 0] OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl ;
 input [ 63: 0] OOOOLL0II0ioIiIIoLOolIOLIoLooIill ;
 input [ 63: 0] OLLI0ilo0LiioOLloOLloiioiIoOiLl0O ;
 input [ 63: 0] OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO ;
 input [ 63: 0] OlOiOoL0i0i0L00OL00l00OOoL0OLILol ;
 input [ 63: 0] OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO ;
 input [ 63: 0] Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l ;
 input [ 31: 0] Ooii00l0ooOoIliILL0lLLLLLoILlIIoO ;
 input [ 31: 0] OILl0LOii0lOi0LlLIIoIL0LLOoli0oll ;
 input [ 31: 0] O0Io0oIliooLo0i0i0lL0IlILOloiiIlI ;
 input [ 31: 0] OLLli0LLl0LlILOoi000iLoiiOOOLooLI ;
 input [ 31: 0] OoIooi0LILolioIilliiol0I0iLoioIoi ;
 input [ 31: 0] OILolilliOIlLILOoioLii0iI0lII0oil ;
 input [ 31: 0] OOIilioOiLLoOIL0iLoILiLLliiio0LOl ;
 input [ 31: 0] OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l ;
 input [ 31: 0] OllioLi0iLLoIOlILoIL0oOO0OiIliOOi ;
 input [ 31: 0] OlOoOLLlO0LOilOiiOoiOi0o0lollolLl ;
 input [ 31: 0] OILoioOioIOL0lIOLoIlIOlolLiOLlIoo ;
 input [ 31: 0] OoI0i0iiiL0ililIOLiL0IioLIL0IooOo ;
 input [ 31: 0] OioIoIoo0iIIlOilLlIoILioo0I0lo00o ;
 input [ 31: 0] OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0 ;
 input [ 31: 0] OLI00Il0O0lI0OoLI0oIloiOIiiILIill ;
 input [ 31: 0] Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL ;
 input [ 31: 0] OioOiiiOlioLLOllo0IiIOiOOli0oi0LI ;
 input [ 31: 0] O0i000LoOoll00lolOOOOIO0Oio0LIO0o ;
 input [ 31: 0] Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO ;
 input [ 31: 0] OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl ;
 input [ 31: 0] Oiio0oo000ioIO0llioIoLILlIlIOOloL ;
 input [ 31: 0] OIooL0lILLIloiOOLiI0ilOIli0LOL000 ;
 input [ 31: 0] OILlOiiL00II0oiOlOoOI0lI00I0oIIIi ;
 input [ 31: 0] OLoOiiL00iolo0LOliOll0I0ILIOL0iLI ;
 input [ 31: 0] OII0Iill0IOLO000li0iL0iLoiIoOoliL ;
 input [ 31: 0] OOI0I0II0oOOO0LiLoO0I00LloOllilIl ;
 input [ 31: 0] OOIioIlLoOL00lOliIIllL00illo0L00o ;
 input [ 31: 0] OLiloooloollOoil0LlolLolOILlO00Ol ;
 input [ 31: 0] OOilLILioilLIliOlOoilOOIolLLiLl0I ;
 input [ 31: 0] OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0 ;
 input [ 31: 0] OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI ;
 input [ 31: 0] OIiLOlOll0ol0OOLIo0oOiIilII0Io00L ;
 input OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI ;
 input Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO ;
 input Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi ;
 input OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI ;
 input OloIioIl0OOlolI0LIiioiLoL0OL0iI0i ;
 input OLIIoil00iiOOl0oloiiooOiI0IlL00Ol ;
 input O0L0oo0LI0OiII0l00oioIIiiilLLIOIl ;
 input OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl ;
 input OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo ;
 input OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI ;
 input OOoo0oiIolLIlol0oll00LiolIOOIlLL0 ;
 input OIlLiI0I0l0olLllLI0LliOOlllliLL0i ;
 input O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o ;
 input OOIILlIiIOiOIi0o0li0lolol0LIoOliI ;
 input OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL ;
 input Ollil0L0OlO0loio0OLiLILo0OioO0iOO ;
 input O0L0O0ioooOOiLLlLLOLiioooILolII0o ;
 input OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl ;
 input OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0 ;
 input OLllIIIO0oIlllOo00LILooILo0io0o00 ;
 input OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI ;
 input O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO ;
 input OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0 ;
 input OllloLIILloiiiOill0lOLooilli0Llii ;
 input OoIL0ll0llIOoI0IoIioiILILllLLOOOL ;
 input OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll ;
 input OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL ;
 input O0oLLI0O0IlOllolLIioIIOll0iiiIlLL ;
 input OiOo0O0ooiioi00lloILL0oLLoILOiLiO ;
 input OlLILiOolLl0ioiLiLlILiILLlIOllloI ;
 input OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O ;
 input O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi ;
 output [255:0] OlolI00LoLoOILILoioLOL0lolLO0oiOo ;
 output [255:0] OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL ;
 output [255:0] O0000Lil0OoOOILlIlOlooioiIOloOioi ;
 output [ 31:0] O00lOOl0oILIoiioLOOI0OoioILioLiiL ;
 output O0iioiILo0ol0ollLilLl0lO0oI0ilOiL ;
 output [255:0] OilO0OLOo0LllI00o0oOil00L0OloIOl0 ;
 output [255:0] OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll ;
 output OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l ;
 output OILLiiO0o00OloIOOl0LlIOOlo00O0OOi ;
 output [255:0] OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil ;
 output [255:0] Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 ;
 output OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl ;
 output Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI ;
 reg [ 1:0] OLILoI0O0oiLILloooL0OLL0iOIoiIoIo ;
 reg [255:0] OlolI00LoLoOILILoioLOL0lolLO0oiOo ;
 reg [255:0] OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL ;
 reg [255:0] O0000Lil0OoOOILlIlOlooioiIOloOioi ;
 reg [ 31:0] O00lOOl0oILIoiioLOOI0OoioILioLiiL ;
 reg O0iioiILo0ol0ollLilLl0lO0oI0ilOiL ;
 reg [255:0] OilO0OLOo0LllI00o0oOil00L0OloIOl0 ;
 reg [255:0] OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO ;
 reg [255:0] OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi ;
 reg [255:0] OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll ;
 reg [255:0] OOollolIl00lOO0iOilIiOol0LOo000iL ;
 reg [255:0] OiILLiLiIiIlIlIOloOlIoOOollIlOiio ;
 reg [255:0] OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil ;
 reg [255:0] OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI ;
 reg [255:0] OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 ;
 reg [255:0] Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 ;
 reg [255:0] Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl ;
 reg [255:0] OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi ;
 reg OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l ;
 reg OioiI0IllllLolOLL0Ii0Oli0lLIL0i0L ;
 reg OLLliiOoIi0oLoIlllooooiLIoLOlL0iO ;
 reg OILLiiO0o00OloIOOl0LlIOOlo00O0OOi ;
 reg OoIoOI0lI0IIIIIoLlOL0o00O0i0OIlio ;
 reg OilL0oiOIollIOIOOO0I0IIoLLOoOOOLO ;
 reg OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl ;
 reg O00oI0oiOi0lLoL0iIL0L0LiLOIlO0O0o ;
 reg OlilIo0olII00llLOlLIloLL0l0iOIOLo ;
 reg Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI ;
 reg O00LIOOl0LOl0OiL0oIOiiOoii00oio0l ;
 reg O0i0oLliiiIoIi0iIi00ILlIooi0OLlil ;
 reg [ 31: 0] OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO ;
 wire [ 31: 0] OiiIlOO0OL0Io00Li00illiLIlIOiLIoI ;
 wire [ 31: 0] Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 ;
 assign Ooli0O0IloLOO0OooL0lIOiiOl000IoO0 = { O0ILIlO0oiLLoOIoIIOliiiilOIlILOoi, OO0IlllIOo0OiilOiOiLI00L0L0OIoI0O, OlLILiOolLl0ioiLiLlILiILLlIOllloI, OiOo0O0ooiioi00lloILL0oLLoILOiLiO, O0oLLI0O0IlOllolLIioIIOll0iiiIlLL, OiIIlLOllOOiIOLIoLOIi0LO00iiOILoL, OiIOiooOOOL0OLoi0ILILlLllLL0l0Lll, OoIL0ll0llIOoI0IoIioiILILllLLOOOL, OllloLIILloiiiOill0lOLooilli0Llii, OLIOIiOL0L0liilOoLLi0lloLiLI0i0L0, O0Lliloi0iIiol0iLIOLlIOOOOOLiOloO, OIlOI0Il0lIlloLoiLolLO0Ll0l0llLlI, OLllIIIO0oIlllOo00LILooILo0io0o00, OO00IIoIiIiIl0IOiIl0oooOI0Lolioo0, OOoi0l0ilLooOII0oIiIlOLO00OOO0oIl, O0L0O0ioooOOiLLlLLOLiioooILolII0o, Ollil0L0OlO0loio0OLiLILo0OioO0iOO, OOoIliLlIoLlo0IlLOIoliioOlOL0o0OL, OOIILlIiIOiOIi0o0li0lolol0LIoOliI, O0iliLIILoiIOlIoO00Ii0OiIoOli0L0o, OIlLiI0I0l0olLllLI0LliOOlllliLL0i, OOoo0oiIolLIlol0oll00LiolIOOIlLL0, OOO00OolOoOlo0OiLi0io0oLoOLOiOLiI, OI0LLOoIOLIOIlIIoLiLOoOIIoiLLLiLo, OoO0LLI0lIiOLL00iOOIooOi0Il0LoIOl, O0L0oo0LI0OiII0l00oioIIiiilLLIOIl, OLIIoil00iiOOl0oloiiooOiI0IlL00Ol, OloIioIl0OOlolI0LIiioiLoL0OL0iI0i, OIoLlOlO0oIoiiLOilooL0IL00LlIiOOI, Ol0OoLIo0IlLlOl0iiOo0LioL0iIllIIi, Ooi0O0iol0IoooL0L00IiOIOiOo0l0OoO, OLoLlI0l0o0iioOI0lL0Ol0IoLOlililI };
 reg O0i0LioOiilLoI00OOLLlio000loo0OIL ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0i0LioOiilLoI00OOLLlio000loo0OIL <= 1'd0 ;
 end
 else if ( O0i00oOl00OoIIOIil0LLOi0looIOIL00|| (|Ooli0O0IloLOO0OooL0lIOiiOl000IoO0) ) begin
 O0i0LioOiilLoI00OOLLlio000loo0OIL <= 1'd1 ;
 end
 else begin
 O0i0LioOiilLoI00OOLLlio000loo0OIL <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO <= 32'd1 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO <= 32'd1 ;
 end
 else if ( O0i0LioOiilLoI00OOLLlio000loo0OIL ) begin
 OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO <= (OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO==32'hffff_ffff) ? 32'd1 : OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO + 32'd1 ;
 end
 end
 assign OiiIlOO0OL0Io00Li00illiLIlIOiLIoI = { OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO[7:0],OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO[15:8],OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO[23:16],OL0ol0oLliLL00OOIiLOlii0oLl0IoLLO[31:24] };
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= 256'd0 ;
 OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l <= 1'd0 ;
 end
 else begin
 OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[ 7:0] ;
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[7:0]) 8'h01: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {OlllLl0L0L0iO0lIloilOOo0iIIiOo00o[23:0] ,OoolLolOioLILoOIII00LIOli00LIlloi[7:0] ,OOOooLlOLO0iOOOLi00oIiloILlooOLIO[31:0] ,OI0lLOI0LIOOil0ioLioLI0OLLliOoI0o[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi[22*8-1:3*8]} ;
 8'h02: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {OOlOIlooi0LiIlLiilOL0LloiII0I0oLo[23:0] ,OOIolooo0Oi00io00lIiiOiiLIliliOio[7:0] ,OlLOO0LloLoiOO0O0i0ilLOi0O00ooiOI[31:0] ,O0oL00IoIIIOLIIlo0oO0lli0ioL00iIi[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi[22*8-1:3*8]} ;
 8'h04: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {O0oLiillllLOiLilOoI000iOLoiL0L0LO[23:0] ,OLLIiolLOOOliIoiIi0oLLiOllooIoiiI[7:0] ,Oo0iOoll0oOLILlOIOI0Oiolol0OlilLi[31:0] ,OO0O0ilLlLII0ilI0oOOOLloilIoOIoLi[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO[22*8-1:3*8]} ;
 8'h08: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {Oio0i0L0iIiIiIl00OIOlOIOlIooIO0OL[23:0] ,OOoL0lOOloLLOLOILLLOolliIll0oOOoO[7:0] ,OIIoiLLooLIIolo0oLiOIoiO0LiiI0lIO[31:0] ,OOllIIoLLLooiiOoLiIi0loOO0ilO00O0[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL[22*8-1:3*8]} ;
 8'h10: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {OoooIiooOl0i0oliO0lio0IOo0iIILLLi[23:0] ,OoOlILlliliiOI0OLLoOOl0000iIo0IIo[7:0] ,OoIlliiIil0Iil00IOL0ooOLIo0O0LiiO[31:0] ,O0lOIi0OI0lOIOIiilL0LOlOIL00oilOO[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI[22*8-1:3*8]} ;
 8'h20: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {OLlLoL0lO0oOIOolIIoiILIO0oOilooll[23:0] ,O0iI0Lil0liLOLiILLOoilII0LII0iolO[7:0] ,OlL0ioloIOIoOLILilIIlIiLo0oIliOLI[31:0] ,OLLIool0I0IooOOIoliL0Oo0iL0L0lOol[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OoIlLi0I0llOlo0lool0LO0O0LlLOILi0[22*8-1:3*8]} ;
 8'h40: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {OiOIlLoIIOoiLL0IOiLIOi0o0LLOo0lIl[23:0] ,O00L00oIOO0IoIOLoLOO0iLiloLi00Lo0[7:0] ,OoLLliL00LLoooll00ooiLolOliOO0lLI[31:0] ,OOLOlIo0lLiLI0I0OLLll0LOlI00io0oi[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OiiOIoolI0LioIo0IlL0lOllILIOOiIio[22*8-1:3*8]} ;
 8'h80: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= {Ooi0Il0iOLOllLLIooO00ilOlo0iOLO0o[23:0] ,O0ooO0I0ii0iiilioiIOO0IlOl0L0lllI[7:0] ,O0li0llLIi0oIo0IilLLooLILolLIOOoo[31:0] ,OioIOIo0IllIo0OILLlli0LOOl00lioII[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l[22*8-1:3*8]} ;
 default: OilO0OLOo0LllI00o0oOil00L0OloIOl0 <= OilO0OLOo0LllI00o0oOil00L0OloIOl0 ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= 256'd0 ;
 OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl <= 1'd0 ;
 end
 else begin
 OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15:8] ;
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15:8]) 8'h01: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {Oio0Oo0Ll0llOOLLloO0LooiiL0LiLOi0[23:0] ,O0II0lLLLo0oiIiiOOLo0OLiOiiiIIIi0[7:0] ,OLoo0OILL0Io0OO0o0oo00OlOOO0LOOOl[31:0] ,O0l0lloOLloIiI0o0LIoi0LOllOIlO0io[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,O0lioOi00lO0IL00IoLLILolIlli00LiI[22*8-1:3*8]} ;
 8'h02: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {OLooLooiioOiOo00LLooO0OLoI0iLiLI0[23:0] ,OIO0IIi0OIooOiLOIII0lLolililiOIll[7:0] ,OioilLoll0OiiOooiLiIOiL0LiilILII0[31:0] ,OLoli0Li0i0oO0olOOilIliIio0LOoIIO[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OOiiIi0oILLIllilLLLOiIi0Ii0lii0II[22*8-1:3*8]} ;
 8'h04: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {Oil0LoiILLliLO0oI0lOIOli0iiOoLOOo[23:0] ,OiLoLLoIoLiooOIIiLOOOIi0oO0oiOiI0[7:0] ,Ol0OLoIiI0OloLIlillLOloLioIIL0III[31:0] ,OiILooool0OiolIOIIlO0LiOliIiIL0Ii[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OoiOoio0IOIoOio0olOLllllOIlLIoiL0[22*8-1:3*8]} ;
 8'h08: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {OLi0ooOo0OlIllLOILllLL00lL00Liii0[23:0] ,OOILOlLi0l0ioiOOIOOI0IlOiiLO0LiLl[7:0] ,Oi0lll0000oiiLo0lOolIi0ooOiiI0lio[31:0] ,OLIIoIiliIoiioIoLoI0LllolIIlO0LOi[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,Oi00i0oL0iIiLll0o0o0l0loi000ioOOL[22*8-1:3*8]} ;
 8'h10: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {OLoI0LiOOoOlLiOLoOI0IOoloL0lLo00I[23:0] ,OO0OOoLL0O0OOOllioILi0liilLLloiLO[7:0] ,OlLlliliOioioOIoiLOIOiOoiiioIOLOO[31:0] ,OIlI0I0IooLOLIlLLLIlli0o0LLl0illI[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo[22*8-1:3*8]} ;
 8'h20: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {OLLoOIOooIOoioOilIIoOlLLOoi0IlI0o[23:0] ,OlL0IOLIoOoilLoIIolLIILoLLI0i0I00[7:0] ,OLoolO0oO0io0IiiiOIIIllllLOO0O0O0[31:0] ,O00IoOolLoIoIoLlIOiOOOoOLl0Iii0O0[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OI0ool0i0ollOOoloL00L0LlLIO0LIliI[22*8-1:3*8]} ;
 8'h40: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {OOIlIio0iILll00lliIIioiIiOLlLLi00[23:0] ,OlIollIiLi0IlLiolloLOOL000Oo0l0II[7:0] ,OIlOoIoi0IoO0iIo0iioLlL0IioILiOLO[31:0] ,OLLiIlIOlII00l00l0LoLLilL0l0OOOLo[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OL0Lio0lIililolilllOL0Li0lIi0I0LI[22*8-1:3*8]} ;
 8'h80: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= {OOiOLoILiiIiOLoOOOl0iOolLLloLLLil[23:0] ,O0oOlLIiOoL0oOoLILI0I0Oll00IlI0OO[7:0] ,OoIIiLoIL0llOo00oIi0oLi00oiill0Ll[31:0] ,OOoLol0oioL0looOlO0io0oIillil0iI0[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0[22*8-1:3*8]} ;
 default: OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil <= OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= 256'd0 ;
 OILLiiO0o00OloIOOl0LlIOOlo00O0OOi <= 1'd0 ;
 end
 else begin
 OILLiiO0o00OloIOOl0LlIOOlo00O0OOi <= |{O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31:24]} ;
 case ({O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31:24]}) 9'h0_01: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OiOO0LOLIOO0LOlloIOIillolO0iIo0I0[23:0] ,OlLIiOlioIILOllO00lLiI0LiIlOloIiI[7:0] ,OllIIoI00oOOiI0LO0OOLiIoiOoOoL00I[31:0] ,OOOOLi0lLIOOoLiioLLoLiLOiiL000OiO[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO[22*8-1:3*8]} ;
 9'h0_02: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OlIli0IolOiL0LoliLloo0olllliIiO0O[23:0] ,OO00il0IO0lLoiilIo0ioiOiOOlLloioL[7:0] ,OLoLOlol00olO0oo0LLlolI0OiLo0llLI[31:0] ,OlIiO0llI0O0Li00OLIILiOLi00OiLioL[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo[22*8-1:3*8]} ;
 9'h0_04: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OIl0iLOOLlOLIIoLLiLilLlLolloIlOi0[23:0] ,OIilIOil0oIoOoo0iiLOIo0L0olo0ooLl[7:0] ,OLolOilolLoloilIloOOiioIloiI0L0Lo[31:0] ,O0lIlL0lLL00000ioioloooIoiiiioi00[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,O0oL00LOlilLooOoiil0oLL0iIillLlLL[22*8-1:3*8]} ;
 9'h0_08: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {Oo0OIlOii0iO0lOIIoli0iOOoLOoOO0I0[23:0] ,O0oIiILIIO0LOOil00IlIoLiIilO00ooI[7:0] ,OiiLlOLO0loioOoLiLIoIiOi0IOIlioLi[31:0] ,OIioLLolLoll0iO0LoLo0ILlii0ilO0o0[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl[22*8-1:3*8]} ;
 9'h0_10: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OoOilOIO0iLL0OLLIo00i0lIlOl0LlOlO[23:0] ,OLOIIIiOOILilol0L0ILiLOiolIl0Oi0l[7:0] ,OO0Oi0ooo0LlLooloL0lLOiiILLi0Oi0o[31:0] ,OioLlLLli0IiOllll0l0LiIoLiLLLOL0L[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OIOio00oLLL0o00LO00LLoI0LlL0OILlO[22*8-1:3*8]} ;
 9'h0_20: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OO00oOlII0oIIIoiOooiIIOlI0Il0l0L0[23:0] ,OoLLOi0lOO0iILIOOliil0o0Lo0IIoLi0[7:0] ,OLololIl0LoiLooLIloiooLli0LOOLLli[31:0] ,OILllI0lillIoilOIoooOll0LII00I0l0[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00[22*8-1:3*8]} ;
 9'h0_40: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OlL0l0OLLIIl0LoLOOLOo0IOiOI0lIoIo[23:0] ,OOIl0oIIIoOLOL00liIiOIo0lo0lIOl00[7:0] ,OIllOIIOiOol000OoLIL0lLl0L00iIIIL[31:0] ,OIIOoooiOOl0l0OlLOlloIlOiI0OOiiLL[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OlLiolooLilLlLiil0l0iiO0IOILool00[22*8-1:3*8]} ;
 9'h0_80: OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {O0lolLi0olIioIiIooOLLLlioIooLIill[23:0] ,OolLO0OOloooOIOiiOilL0IiILL0iol0I[7:0] ,OL0looio0Loioi0ill0olOo0o00ioOOII[31:0] ,Oo0o0ooIOoiiLIoloLoLOoOOliLoiO0OI[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i[22*8-1:3*8]} ;
 9'h1_00 : OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= {OLO0oOILL0O0IIOOiLlLOoioI0iiiOOiI[23:0] ,OilIL0OIOillLolooIl0LLIo0lIL0Ooo0[7:0] ,OLoIlIiLIIIoI0oIOillIIOOLoIIoO0ol[31:0] ,OloliIooiiLI0IIlOiL0LLlioILLllL0L[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OioILlIiO0000OoolooO00loIOIloLIoI[22*8-1:3*8]} ;
 default : OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll <= OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= 256'd0 ;
 Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI <= 1'd0 ;
 end
 else begin
 Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23:16] ;
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23:16]) 8'h01: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OLio000LoL0lOol0oIiLlILLIlOLLOIlO[23:0] ,OOoIIOoIl0LIOllIO0L0oLoOIOoooiill[7:0] ,OIO0l0IOIol0iIl0i0oiliOioLLLi0Ili[31:0] ,OILIi00LOILOoLIiLloLiLIolliOoooIo[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OI0L0iIOilOi0LlILL0l0liiiil0lOIii[22*8-1:3*8]} ;
 8'h02: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OoiiooOo00OI0O0loiolLOLioIOiI0LoI[23:0] ,OiOIOlILOi0lIoOiIOIoOIllLILLiIliL[7:0] ,O0IIL0iIliIIolLLiioLIILlIoI0o0IOI[31:0] ,OIi0liIIIoiOooLllLO0O0IoLLllIOlli[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL[22*8-1:3*8]} ;
 8'h04: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {Ol0L0iLLLLLLLo0IlIoI0liLLIiolilOl[23:0] ,OO0LO0iliiL0Oi0OIIloILLOiO0LLloli[7:0] ,O0ilOlIii0IliiO0OoiIi0oLol0L0lLiO[31:0] ,O0ioIo0IOoIIOOlIIOo0l000LI0iio0iI[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OooOIi00Ii0liOollOoLioI0OiLiLiO0O[22*8-1:3*8]} ;
 8'h08: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OOLooiiL0oLlI0Lo0I0LiL0o00LllLO0I[23:0] ,O00OiooIolIi0oIoIiiLlO0IiIO0ooLio[7:0] ,OO0llOooLooLoi0l0oIOOoilOolIoLLOo[31:0] ,OOIIlilOoOlIolLlILLioil0LL0oLlloo[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol[22*8-1:3*8]} ;
 8'h10: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OIO0IioIOoIOIll0LOIlOOILoILoiilli[23:0] ,Oo0i0IlILOo0ooOiIlLOoiioll0LilllO[7:0] ,OLl0oiiIOL0ol00LIoo0IoolIollol0ii[31:0] ,OLiiOLILl0LIlL00OlL0Oili00IiIlIl0[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OiILIII00lOolOiililIOiIIloo0OlLlo[22*8-1:3*8]} ;
 8'h20: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OLoOLiILLLiIilOolo0Lil0iLLOOLILII[23:0] ,O00liliooOOoiI0OlOOIIlO0o0IiOOolL[7:0] ,OILLl0iillioLoOiiIiL0iliIOiO0oiio[31:0] ,OOLOoOLoILILOOL0OLL0i0lLI0Oi0LlIL[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OiioOooilOllI0oOoolilo0OLIlioo0II[22*8-1:3*8]} ;
 8'h40: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OOoLoi0LlLLLoIIllLLLIli0OI0LlliII[23:0] ,O0IOLlLLoiioi0LIOo00oLLOlOLL0oooI[7:0] ,OIIOOOiLO0IO0I0oIIOolIOLlLOLi0oI0[31:0] ,OOiOiIiiilililLoLlIOoIoiILilLoooI[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OIiolOOI00iliL0LolLOOOLOliiIlLlII[22*8-1:3*8]} ;
 8'h80: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= {OiLl00LLioIio0iLiOiIOOOlLIlilOIOi[23:0] ,Oil0LOOoLO0iIOooiIiO0IlilOLIlIoOO[7:0] ,OOoILooiOiiiIll0oOLLIIoO0oLolIIo0[31:0] ,OO0O00OIoioOIOLi0IlILI0OlilooOIOo[7:0] ,OiiIlOO0OL0Io00Li00illiLIlIOiLIoI[31:0] ,OLOL0OioiLOLoli0LOL00OOiO0iiOooll[22*8-1:3*8]} ;
 default: Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 <= Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlolI00LoLoOILILoioLOL0lolLO0oiOo <= 256'd0 ;
 end
 else if ( OiiIOOL0iLil0OIO0OLlOiLiIOolO0i0l ) begin
 OlolI00LoLoOILILoioLOL0lolLO0oiOo <= OilO0OLOo0LllI00o0oOil00L0OloIOl0 ;
 end
 else if ( OILLiiO0o00OloIOOl0LlIOOlo00O0OOi ) begin
 OlolI00LoLoOILILoioLOL0lolLO0oiOo <= OOiLLOl0lIoOiL0IIOl0lOoIlilIiI0Ll ;
 end
 else if ( OiIil0Ll0lIlOlillOLiLOoOoiIlO0IIl ) begin
 OlolI00LoLoOILILoioLOL0lolLO0oiOo <= OOOl0LIiLolLiiLiIlIoIlIioIOLIiOil ;
 end
 else if ( Oiilioi0OOo0LI0I0LOi0OOlLI0IOIooI ) begin
 OlolI00LoLoOILILoioLOL0lolLO0oiOo <= Oo0IooOlLiiL0oIll0LIoo0iOlL0LO0i0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= 256'd0 ;
 OioiI0IllllLolOLL0Ii0Oli0lLIL0i0L <= 1'd0 ;
 end
 else begin
 OioiI0IllllLolOLL0Ii0Oli0lLIL0i0L <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[7:0] ;
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[7:0]) 8'h01: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {Oll00l0Lo0l0iLLLOIOLoL0io0OLLLooi[3*8-1:0] ,OLlIOIOlOLllLii0IoI0oiOIOiiLoiOI0[71:0] ,OIiO0OLioLiIOIIiLoiLooI00I0olI00O[31:0] ,OOOo0I0LlloiIl0i0il0OLiOlooOOolil[63:0] ,OO0LLiOLIi0liI0LolIoLiIolOoi0Ii0o[31:0] ,OLlOlii00IoIl00oIioIiIool0lLiOoLo[8*8-1:4*8] } ;
 8'h02: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OOIliLOooOOIoIOOOllLiIIlI00Ol0iIi[3*8-1:0] ,Oo000ooL0O00L0illOlOLOO0oilOIi0Ll[71:0] ,O0Ol0i0loLlooOIiLoOlIilLolOlio0ll[31:0] ,OoiIO0i0oolLLiLllI0OI0lio0Lo0i0Li[63:0] ,OoI00LooIIlIIlIOOLIoloilI0OoIILLi[31:0] ,OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL[8*8-1:4*8] } ;
 8'h04: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OiolOoioIIl0ILO0OIOoIOioOiiOoiIOO[3*8-1:0] ,OlIloooO00OIL0L0iIili0iOOoiLI0oiI[71:0] ,OOIOoLoIIIiiLLOLIOloiLIOi00oi0L0I[31:0] ,OolIilIL0iooOLllOLloloOIlLIiOoLo0[63:0] ,OIoIo0LOLLil00oOL0ILoI0OlOOiLOLII[31:0] ,OL0LLioOOooILOL0LLLIilLl0oLLiIoiL[8*8-1:4*8] } ;
 8'h08: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OOiLilOOiIOLL00OlOi0OLlL0ioIIOoIL[3*8-1:0] ,O0OLLIlOIIi0iL0ioIiooOOil0ILo0LIL[71:0] ,O0ioIlLL0lloioL0LoiLoLLloL0OI0ILi[31:0] ,OOOLoOoloOlLiL0l0IIOolOlioLLo0LlO[63:0] ,OL0OIiOoo0IllO0oloolIll0oOo0LlIIi[31:0] ,Ol000OloII0LlIII00IIOIlOiioOo0Iii[8*8-1:4*8] } ;
 8'h10: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OLiIo0lIo0iOLiOiiO0L0lOo0OooIL0LI[3*8-1:0] ,OLolLol0lLIIlIillI000oIlilLLloOii[71:0] ,OiOiOiIIiLi0OIILO0Ioi0iLl0ILLOOoo[31:0] ,OoIiLlLoiLlOl0oLOlIIoO0l0lIILLI00[63:0] ,OO0O0oOlliIoIOlooIO0lOLolIilLllIO[31:0] ,O00I0iOoILll0oILl0ILloii0LIIOOiIO[8*8-1:4*8] } ;
 8'h20: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OoIlLi0I0llOlo0lool0LO0O0LlLOILi0[3*8-1:0] ,OoIoIO0O0oOoilLlI000OIllIIoI0ioIl[71:0] ,OLLloO00IliLiLLlLloLloO0liOoIIOOI[31:0] ,OooL0L0LLLOoL0IooiiiO0OLOIiiO0OLl[63:0] ,OOIlLIiol0o00OlI0lLl0lILiIolL0iIi[31:0] ,OO00IIiOlOioiOLIiIloilLII0lLL0OOi[8*8-1:4*8] } ;
 8'h40: OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OiiOIoolI0LioIo0IlL0lOllILIOOiIio[3*8-1:0] ,OoIooolIllLIIolLII0IiLLiiOlOOIIOO[71:0] ,OL0OIO0I0IOoOoiIOllLIOlO0lio00IOi[31:0] ,OLL0i00LllLlio0oLOLooIL0ilLLllil0[63:0] ,OOiOiOIIoOii0oOLlI0OliIi0liioLLII[31:0] ,OlOl0iOIioolOiill0OLOloOoLiIlllol[8*8-1:4*8] } ;
 8'h80 : OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= {OlL0O0OiOIiilOOIooIlo0lO0li0oOL0l[3*8-1:0] ,Oli0oLliOoIo0IOoIOiLLIlIioLiIlLio[71:0] ,OOI0o0iiIlloiiIoiolooi0Ii0IL0oLOI[31:0] ,OLLLllOIlLOioiIIoOIOiLOILOioLlLLo[63:0] ,O0oiILoiiI0oOOoiillLOoiIilI0o0Ool[31:0] ,OOooOoIiooIliiO0LoLiOlOoIlOOo00I0[8*8-1:4*8] } ;
 default : OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO <= OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= 256'd0 ;
 O00oI0oiOi0lLoL0iIL0L0LiLOIlO0O0o <= 1'd0 ;
 end
 else begin
 O00oI0oiOi0lLoL0iIL0L0LiLOIlO0O0o <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15:8] ;
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15:8]) 8'h01: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {O0lioOi00lO0IL00IoLLILolIlli00LiI[3*8-1:0] ,OI0i0lOolo0oOILo00ll0LIIOiOOlIoii[71:0] ,OOiiolOoloIoil0iO0OiOIIoL0OlO0o0L[31:0] ,OL0oloO0o0o0oli0I0IOo0olOLLoLOl0I[63:0] ,OI0O0lOIO0OOOOllIL00Ooi0I0llLlili[31:0] ,OioOlIooLl0IL0LiioIlILIolO0o0ii0l[8*8-1:4*8] } ;
 8'h02: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {OOiiIi0oILLIllilLLLOiIi0Ii0lii0II[3*8-1:0] ,OIILOOOOIOl00OoIollioiiliIilolLLl[71:0] ,OiooooLLoI0OLilIIil0ilooLo0OIloLl[31:0] ,O0iooIILOi0llLIIoILoo0ilIIIlooLI0[63:0] ,OiLiiLILIoLilioiLolliOl0LI00LLil0[31:0] ,Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0[8*8-1:4*8] } ;
 8'h04: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {OoiOoio0IOIoOio0olOLllllOIlLIoiL0[3*8-1:0] ,OO0OIIllLILi0iIlOOoLIIiOoL0oolOL0[71:0] ,OIoLIIo0iOIloioO0IlLoOOliLoIoI0LO[31:0] ,OlI0L0O00L0O0oIIlioOl0ioOIoiIoIL0[63:0] ,OLlolloLliiLO0IlIlLo0lIiiloL00OOL[31:0] ,OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO[8*8-1:4*8] } ;
 8'h08: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {Oi00i0oL0iIiLll0o0o0l0loi000ioOOL[3*8-1:0] ,OOIoiLiIoOOiOIIoLOliOLO00i0IoII0L[71:0] ,OOOLilOolI0LILLIoloIiO00OiIiLiiIo[31:0] ,OIoLOOIo0i0iLiOiIIO0II0LIiiiioIOl[63:0] ,OooLI0lioLIOiOOI00oLLOiLIOlO00ILi[31:0] ,OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol[8*8-1:4*8] } ;
 8'h10: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {OoLoilLlI0lOIOliOl0I0lLOLLLiLILoo[3*8-1:0] ,OooiL0oOLIIOoi0liOLiLOiLIOIILLo0L[71:0] ,OolOi0LliLO0iiLI0oLIlilIlIIIOlL0l[31:0] ,OliliILl0LLiioool00L00LoLLILio0lO[63:0] ,OL0Oloi0OoLOiO00LLloIolIo0iiLLOII[31:0] ,OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII[8*8-1:4*8] } ;
 8'h20: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {OI0ool0i0ollOOoloL00L0LlLIO0LIliI[3*8-1:0] ,Oo0loliLllliloIiliOi0lILloLI0ILlO[71:0] ,Ooi0OL0i0IioliooLiI00OoiL00looOIL[31:0] ,OliiIiOLlOL0Ii0IOioIIoIL0ILo0OL0O[63:0] ,OOo0lLI0lLOLIOILoo0I0o0iOLIILoiIo[31:0] ,OoLO0LoiiIL0lilol0oloO0loiLLiIIl0[8*8-1:4*8] } ;
 8'h40: OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {OL0Lio0lIililolilllOL0Li0lIi0I0LI[3*8-1:0] ,O0OI0iLlL0LOLlOolLOoLLILLoI0lo0io[71:0] ,OolL0oo00LOo0LOoLiILllLo0loOoIiii[31:0] ,OIOIOlilIolIlLOLlLlll0IiOIiILiOol[63:0] ,OiloLLIlO00Il0oo0io0Iilliiil0OolO[31:0] ,O0oOL0illOloooo0ioIiOLOooLILllLl0[8*8-1:4*8] } ;
 8'h80 : OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= {OIlIlo0IO0LIIoO0LlLOLOloOIL0OlLL0[3*8-1:0] ,O0oilLoOiOiLLi0Li0lLOIooIiliILlii[71:0] ,O0o0OLOoLlLiL0oiI0Li0lOoLO0LlOi0l[31:0] ,OL0Ool00li0LiiLlOiOooIOi0i0LOlIoo[63:0] ,OLI0iO0OLLO00l00LIlOLiiLlloILOLIl[31:0] ,OLiILioillIololIOILoOLlI0LILLliIL[8*8-1:4*8] } ;
 default : OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI <= OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOollolIl00lOO0iOilIiOol0LOo000iL <= 256'd0 ;
 OoIoOI0lI0IIIIIoLlOL0o00O0i0OIlio <= 1'd0 ;
 end
 else begin
 OoIoOI0lI0IIIIIoLlOL0o00O0i0OIlio <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23:16] ;
 case (Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23:16]) 8'h01: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OI0L0iIOilOi0LlILL0l0liiiil0lOIii[3*8-1:0] ,OlIIioIIlILoli0oIiIl0l0IlOlloooll[71:0] ,O0LiloL0oiioIoLlOLlIIiiIOOl0Lli0I[31:0] ,OO0loiO0lOooolLIoOIoOLlOoLlO0ioL0[63:0] ,OLIOiIoLIlIo0liLIOii0ilLiiiIOL00I[31:0] ,Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0[8*8-1:4*8] } ;
 8'h02: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OIlIlO0oiLILoIIoLlIoioI0II0iL0LOL[3*8-1:0] ,OOL0LIooi0LlIli0I0ooO0LiOI0IIliOO[71:0] ,OllLlOiLLooiILOiiOOlLlL0LOII0LLOL[31:0] ,OI0OLOILiOlOoolLIilooolollLLo0OOO[63:0] ,O0Il0L0lLloiIiliL0000o0oIOLLILool[31:0] ,OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0[8*8-1:4*8] } ;
 8'h04: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OooOIi00Ii0liOollOoLioI0OiLiLiO0O[3*8-1:0] ,OioolLOlII0IlolOIiLOliilL0oiiOoIo[71:0] ,OilO0i0Lll00Iolo00lOOLiLiOiLO0lio[31:0] ,OoII0il0iLlL00iIo0I0OoloiiilLOLIo[63:0] ,OiI0ILIIIiiLO0LOlOLliioLL0II0OooL[31:0] ,Oi0Liloll0L00OiL0iLli0LO00iloIoLi[8*8-1:4*8] } ;
 8'h08: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OilllIOiIlOoIl0oOLOiIOlOOlLi0I0Ol[3*8-1:0] ,OLIoilIIoI0Ol0Oll0I0LloliiLlolIII[71:0] ,OILi0IiLoLOllLioi0oiOlIILl0oiOoi0[31:0] ,Ol0L0l0iLL0LiOOIL0oI0OOolLoiOli0l[63:0] ,OOoooLL0l0llOLI0o0oO00LIoLO00LILO[31:0] ,OoilLIlliloO0LoOL00IILioiolLIloi0[8*8-1:4*8] } ;
 8'h10: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OiILIII00lOolOiililIOiIIloo0OlLlo[3*8-1:0] ,OL0IOILllOOO0OIOL0000LoO0llOo0Lo0[71:0] ,OLOl00iiILoiI00i0lOlLOi00IOLLlOIL[31:0] ,OIooL0i0o0o0OlIioiil0lOoIiI0OLlOl[63:0] ,OioIOlLLLIoiIilLOoiIOIOI0ilI0ILLl[31:0] ,OLIloIl0iIiooOIo0lLlO0L00LOIil0LO[8*8-1:4*8] } ;
 8'h20: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OiioOooilOllI0oOoolilo0OLIlioo0II[3*8-1:0] ,OIolOIIiLIloloOL0iIIO0il0li00ilOo[71:0] ,OlOllIloiIIIIloliooOo0LoIil0o0oii[31:0] ,OLIoLi0ioO0OLLl0LlIOillIoili0OIOI[63:0] ,OIIooiOIlLOiLooO0ioOiIiILOiLLO0L0[31:0] ,OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO[8*8-1:4*8] } ;
 8'h40: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OIiolOOI00iliL0LolLOOOLOliiIlLlII[3*8-1:0] ,O0lIoLOO0iiooiliLlIoiloOLOlLO0IiO[71:0] ,O0OoiooiIOLOllil0OLoLOlllL000LII0[31:0] ,Oi0oIIOolOLiiO0OI000OLlI0OOiIlo0i[63:0] ,OOl0i0OIIooLiI0IioL0LLILIloOlOllL[31:0] ,OOOlLolILloIii0oollOil0lI0OOoOoo0[8*8-1:4*8] } ;
 8'h80: OOollolIl00lOO0iOilIiOol0LOo000iL <= {OLOL0OioiLOLoli0LOL00OOiO0iiOooll[3*8-1:0] ,OILl0Ol0LliiIi0IlOlO0llOlliLlOo0L[71:0] ,O0oiOOLLiiillOliOOOllO0iO000OOoLI[31:0] ,OIliOOilOillIo00oiOOLIOiLolIIooOl[63:0] ,OIi0IoOiOolIo0LlLLOILoLlIliIiOOOO[31:0] ,OIlOIiiliIlIOIlilliilOl0iILIOOOLO[8*8-1:4*8] } ;
 default : OOollolIl00lOO0iOilIiOol0LOo000iL <= OOollolIl00lOO0iOilIiOol0LOo000iL ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= 256'd0 ;
 O00LIOOl0LOl0OiL0oIOiiOoii00oio0l <= 1'd0 ;
 end
 else begin
 O00LIOOl0LOl0OiL0oIOiiOoii00oio0l <= |{O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31:24]} ;
 case ({O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31:24]}) 9'h0_01: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {O0oIoIlILoII0Oi0i0lO0oLLoil0l00lO[3*8-1:0] ,OOIIOLL0llI0lLoloO0ioL0OLLOLi0ILl[71:0] ,OlIIloOL0iLIOLlOlLILlloiioloooILi[31:0] ,OolOOLl0OlII0OiiloIloOO00IllliiLO[63:0] ,O0oIOOiI0OiOlLoo0o0oiloL0oIiOIo0O[31:0] ,OIliolloLooOi0OolOOi0ILOlIliLi0o0[8*8-1:4*8] } ;
 9'h0_02: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {OiI0iO0oL00oIolOOoLOiI0I0lOoilLOo[3*8-1:0] ,OLiLLLlIIIII0LI0LloIIOLi0LlOioIIL[71:0] ,OOLLIiOOi0IloO0I0Lo0oOiillLIOol0l[31:0] ,O0o0OillO0LllooIiILLoilol0lii0liL[63:0] ,OIO0L0iO0iLllOLILO0IoLliLolI00lLI[31:0] ,OI00OOL0LLOOLLLiIooi0oL0iioOloL0O[8*8-1:4*8] } ;
 9'h0_04: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {O0oL00LOlilLooOoiil0oLL0iIillLlLL[3*8-1:0] ,OoILi0Ii0lllOoioI0Ii00LIOLoOIo00L[71:0] ,OOILlooOIliLloiliIOi00LIlLIoli000[31:0] ,OLOlILilLoI0liOiooL00OOlo0i0LiiiI[63:0] ,O0oOLILIoIlLOIIollLOoL00o0O00OiOo[31:0] ,O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L[8*8-1:4*8] } ;
 9'h0_08: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {Oio0lo0iLOiilILL0IlIoi0OIoi0LLLLl[3*8-1:0] ,OIL0OiIiiiOLliIioloLo0lLILolLoLL0[71:0] ,OiIL00IOiOiiI00oiio0lLOlooIiLiOio[31:0] ,OOIIilloi0OiOoo0iI0LI0LI00oILiLio[63:0] ,Oi0OlLiOoOoLLOiolOIOllIoo0LloOIIl[31:0] ,OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0[8*8-1:4*8] } ;
 9'h0_10: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {OIOio00oLLL0o00LO00LLoI0LlL0OILlO[3*8-1:0] ,OILLLoLI0LiOLilloOiLOIlILI0Io0l0o[71:0] ,O0iIoLOl0iLLIlIoOLIol00OlOiol0LIo[31:0] ,OI00OlliiO0LlIIiOoIL0oooi0LloLLo0[63:0] ,OoooO0olOolLIIOLIIl0L0ooLIOoOOioL[31:0] ,O0illollo0oliIl0OolOoIlIILL0OIioO[8*8-1:4*8] } ;
 9'h0_20: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {OlLiOLlii0Oi0LLliLlL0OLioILi0Oi00[3*8-1:0] ,OoII0IlLLoIio00Ii0iOlLIOLIiiL0LIl[71:0] ,OilIl00OOIloIli0LIIii00LIIlILiL0L[31:0] ,OOLiOLLli0OOIOOIo0l0O0O0I00l0LO0O[63:0] ,OOl0LLoL0ioo0iLILI0i0ooLLL0io0l0o[31:0] ,OoOoIOoI0LILoIlIliLIioOooOOOIOoli[8*8-1:4*8] } ;
 9'h0_40: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {OlLiolooLilLlLiil0l0iiO0IOILool00[3*8-1:0] ,OoI0I0oILOoOo0OOIOl0LIolOiOl00IoI[71:0] ,OLlO0iOoIoLLOOii00OO0iLo0oIlOo00I[31:0] ,OIoolOll00LlI00l0oIOLLIOI0I0LIILo[63:0] ,OliiLIIoII0Lo00iio0O0iiIlI0ooIiI0[31:0] ,OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L[8*8-1:4*8] } ;
 9'h0_80: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {Ol0o0OiIIII0iIiiIOOoIIo0llolIoo0i[3*8-1:0] ,OI0oL0loOli0oOIo0oi0lLlolOOiooIo0[71:0] ,OO0oIOllioLiLlLLlii0ilL0OlIliIilO[31:0] ,OlO0LlOLl00IIOIOiilooOLo0liLiIOl0[63:0] ,OLoOO0OOIooLoI0liLOLllIiIOIL0Olol[31:0] ,OLOllOoI0IolOloolLolO0lIiolLiIILi[8*8-1:4*8] } ;
 9'h1_00: Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= {OioILlIiO0000OoolooO00loIOIloLIoI[3*8-1:0] ,OLOl0000OLooLIIo0lIOIOI0lILioolOl[71:0] ,OIiL0oOlOl0iOLIiilOol0oIoOL0L0iII[31:0] ,OoIolLlOIIoIoi00lloLlIoI0lo0iILol[63:0] ,OLiILI00I0Ii0LolLL0oLoLl0IIolOOiI[31:0] ,OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[8*8-1:4*8] } ;
 default : Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl <= Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL <= 256'd0 ;
 end
 else if ( OioiI0IllllLolOLL0Ii0Oli0lLIL0i0L ) begin
 OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL <= OlO0oOOiLLOoLlOi0Iolo00LLoiIOlLlO ;
 end
 else if ( OoIoOI0lI0IIIIIoLlOL0o00O0i0OIlio ) begin
 OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL <= OOollolIl00lOO0iOilIiOol0LOo000iL ;
 end
 else if ( O00oI0oiOi0lLoL0iIL0L0LiLOIlO0O0o ) begin
 OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL <= OOli0iLOIOIoIi0ilOl0oiLOI00OIO0lI ;
 end
 else if ( O00LIOOl0LOl0OiL0oIOiiOoii00oio0l ) begin
 OlLL00ILioO0IiO0OIOI0oolLL0IiLLiL <= Oloi000LiLlIl0iO0LIIllOiLOoOIOIIl ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= 256'd0 ;
 OilL0oiOIollIOIOOO0I0IIoLLOoOOOLO <= 1'd0 ;
 end
 else begin
 OilL0oiOIollIOIOOO0I0IIoLLOoOOOLO <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23:16] ;
 case ( Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[23:16] ) 8'h01: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {Oo0lIOlIlloLIo0lLooL0liI0lIIiLLl0[4*8-1:0] ,OIOO0oiiIiiOILOOioiiO00OIl0lilllO[8*8-1:0] ,OOLlI0LIiLl00iLol0oLiiOoOiiiOIloO[8*8-1:0] ,OO0iLILOLioOioLOoLIOlOlo0oOIollll[31:0] ,OI00OlLIOIiOOiIliIooII00LLLllLLOO[63:0] } ;
 8'h02: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {OOOIioIlO0LIlL0llOIOIOIL00IOIoIi0[4*8-1:0] ,Oo00IIIIoOIO0IL00llOoOioiollIOi00[8*8-1:0] ,OlIliOioiio0LLoLl00i0liioIOI00iIi[8*8-1:0] ,OLOlLlooLIlL0IIiOilIiIooLloIioLOi[31:0] ,OOlOiiLoIooll0L00oIIIoOIililiillo[63:0] } ;
 8'h04: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {Oi0Liloll0L00OiL0iLli0LO00iloIoLi[4*8-1:0] ,OolIl0OOoiOlLioiloO0OolLOiIOolLLI[8*8-1:0] ,OOiiILOoLlI00LoOil0OiOoIlloIiOi0o[8*8-1:0] ,OOl0oiloLLLIo0Li0ioloOiioLl0I00O0[31:0] ,OlIOlLIlLOIlLio00OIiLloIooIOo0ol0[63:0] } ;
 8'h08: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {OoilLIlliloO0LoOL00IILioiolLIloi0[4*8-1:0] ,OL00oOoLi0iLl00LILOOLOlooiiLOOoLo[8*8-1:0] ,O0ioLLo0liLOOiOL0OoLiOool0lLI00oi[8*8-1:0] ,OoIlL0lI0iL0iiIoLii0lLLio00lIIOol[31:0] ,Oll00iO0Ol0IOLloLLilo0OliIloIiLli[63:0] } ;
 8'h10: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {OLIloIl0iIiooOIo0lLlO0L00LOIil0LO[4*8-1:0] ,O0lIi00lIl0iOlLilOloOIllllLLolooo[8*8-1:0] ,OI0O0oLO0looiLoLIL0ii0oIOlI0Lo00o[8*8-1:0] ,O0O0L0iLLIlOILiOLoIiLiliiIllIi0li[31:0] ,OIl0iolIOLOlLOloIoLoIo0OooLi000lO[63:0] } ;
 8'h20: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {OilLiLlOlOLLlLlil0IIiiLiiLlILlIoO[4*8-1:0] ,OoO0ooI0oo0OO0lioOLLlol0L0iOi0OOL[8*8-1:0] ,OLILoOooIiil0oIIolILIlLIioL0i0Iio[8*8-1:0] ,OOLIlOoI0oOlII0oIllLi0l00iOioLIOi[31:0] ,OoiIOl0lloi0IiIlIILIIIIOLloL0LLlI[63:0] } ;
 8'h40: OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {OOOlLolILloIii0oollOil0lI0OOoOoo0[4*8-1:0] ,O0IOiLlL0I00Iol0LiLIOoILiLII0LiI0[8*8-1:0] ,O0lLOioIo0oiOLiollIOLioI0Ii0iLi0O[8*8-1:0] ,OOI0llLoO0IOO000OilllLLLI0i0Iilil[31:0] ,OOIOl00lliliioILLoiioolL0OLLoLo0i[63:0] } ;
 8'h80 : OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= {OIlOIiiliIlIOIlilliilOl0iILIOOOLO[4*8-1:0] ,OIoll0OLiliiLlIililii0oiII0Ol00lO[8*8-1:0] ,Ol0LliIIIIiOOILo0ooioLolOOOololIo[8*8-1:0] ,OlollLLLoL0iiI0lool0OOOOIiOoolioL[31:0] ,O0LLLIIil0l0lOIo0llOLo0oOI0iiIIL0[63:0] } ;
 default : OiILLiLiIiIlIlIOloOlIoOOollIlOiio <= OiILLiLiIiIlIlIOloOlIoOOollIlOiio ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= 256'd0 ;
 O0i0oLliiiIoIi0iIi00ILlIooi0OLlil <= 1'd0 ;
 end
 else begin
 O0i0oLliiiIoIi0iIi00ILlIooi0OLlil <= |{O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31:24]} ;
 case ({O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[31:24]}) 9'h0_01: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OIliolloLooOi0OolOOi0ILOlIliLi0o0[4*8-1:0] ,Ol0IO0lOlO0O0lilIOLiO0L0lilio0LOi[8*8-1:0] ,OIILiOiLOO0IILI0llIOoooi0oLiiOioO[8*8-1:0] ,OLOILIii00lILOLoLIIlOiioll0ilOLii[31:0] ,O0IlliiI0l00iOLL0oLilIILo00lLIolo[63:0] } ;
 9'h0_02: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OI00OOL0LLOOLLLiIooi0oL0iioOloL0O[4*8-1:0] ,OoOll0iOi0l0LiioLllOoliOoO00Lloil[8*8-1:0] ,OiIoioILioOLl0io00oiOiO0liliOlOoO[8*8-1:0] ,OoLI00lolL0IOil0OOLOOooLLIIOOl0Ol[31:0] ,OIioI0IoIoL0ILiiOIOoiO0OOliIIoiOl[63:0] } ;
 9'h0_04: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {O0I00lliIoIlOLIolIIi0ooiLlO0l0L0L[4*8-1:0] ,OOIoI00iO0IiilOOoILo0O0O0Oioo0oO0[8*8-1:0] ,O0OOOLLL0oOLoillIiOLIiIoI00LioiLl[8*8-1:0] ,O0OllOiIO00LliIOoLolo0loIiL0LiIlI[31:0] ,OOOOLL0II0ioIiIIoLOolIOLIoLooIill[63:0] } ;
 9'h0_08: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OlLo0IiIiliLoI0O0lIoliOLLO0ILL0O0[4*8-1:0] ,O00o0iOOoOiLI0iiIOoIiIliLoIliIIll[8*8-1:0] ,Ol0lLoOLiiLllLOoL0OI0Iil0OloOLlLo[8*8-1:0] ,Ooo00lolOl0OIoLOIlIliL0oLooIolLiL[31:0] ,OLLI0ilo0LiioOLloOLloiioiIoOiLl0O[63:0] } ;
 9'h0_10: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {O0illollo0oliIl0OolOoIlIILL0OIioO[4*8-1:0] ,O0Il00oIILloI0IL0LiOO0i0lIiIoolio[8*8-1:0] ,OiLlO0oiOoiLoIIlOlIoOoO0l0OLO0loO[8*8-1:0] ,OLoiiLOLoLOl0lO0LIL00OIolLIo0iOol[31:0] ,OIlo0IlilLOloLLiLIiOOILOLOIl0LOIO[63:0] } ;
 9'h0_20: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OoOoIOoI0LILoIlIliLIioOooOOOIOoli[4*8-1:0] ,OI00OLIIi0LioLLLLllooOiOl0iolOO0I[8*8-1:0] ,OiilOlIoIIlLL0l0I0IlIIIO00O0oliiO[8*8-1:0] ,OLIIl0o0liIOIooiOII0liO0oLllOI0oO[31:0] ,OlOiOoL0i0i0L00OL00l00OOoL0OLILol[63:0] } ;
 9'h0_40: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OiOIoLOiiLOl0oil0IILLIi0IIoLlLI0L[4*8-1:0] ,OO0IOiiiiOIlLLIlIOLlOlII0iiLlOliO[8*8-1:0] ,OLilli0Oo0Ill0lIoO0oILoLLiioOiLiO[8*8-1:0] ,Olo0llLLi0L0IiLooLi0IooLOol0iIiIO[31:0] ,OOLOoLoLOiOOOILIiOoOOLiOLOlLoIOiO[63:0] } ;
 9'h0_80: OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OLOllOoI0IolOloolLolO0lIiolLiIILi[4*8-1:0] ,OOILLooOOlllIILoIiIioLIOI0LOiLiLI[8*8-1:0] ,O0iOioiLIOo0OIloIlIi0OIoO0i0ILIIi[8*8-1:0] ,OOo0ollLl0iLoOI0liLlOoLoL0OLi0i0O[31:0] ,Oo00oLIOoIlL0ooIOIoooiolO0oIOOO0l[63:0] } ;
 9'h1_00 : OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= {OlolLoOiilOi0I0I0I0I00L0LIIILI0Lo[4*8-1:0] ,OOIIloOlOILliIOILOIOiIlooIOOIL0oO[8*8-1:0] ,OllLi0iLIIoo0LOioloOlIO0IlOO0i0Io[8*8-1:0] ,OiLOo0loOI00OL0Ooio0OIIlOLiooLOII[31:0] ,OlLilll0ilOLI0IIoO0li0l0OlO00oLIO[63:0] } ;
 default : OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi <= OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= 256'd0 ;
 OLLliiOoIi0oLoIlllooooiLIoLOlL0iO <= 1'd0 ;
 end
 else begin
 OLLliiOoIi0oLoIlllooooiLIoLOlL0iO <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[7:0] ;
 case ( Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[7:0]) 8'h01: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {OLlOlii00IoIl00oIioIiIool0lLiOoLo[4*8-1:0] ,OIollo0oLlLiI0IILOO00illIILLIoo0o[8*8-1:0] ,O0Lo00iLoOIlILilLooLoiOLi0ooi0iOL[8*8-1:0] ,OIOIIiIlOo00OLl0lOL0IiLOloLL0OOoi[31:0] ,OLli0lIO0lOO0OooILllIi00Lol00oili[63:0] } ;
 8'h02: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {OL0oLOoLiiIioOOiLLLOliL0o0LOIoolL[4*8-1:0] ,O0LIlOOoIoIllLoI0oooOiLoOoIlILLi0[8*8-1:0] ,OOIoOIilLi0looLILloOOollIIIo0llLo[8*8-1:0] ,OiLiOiL00IOIl0loOiOOOiOIlllIOL0iL[31:0] ,OOllI0oo0L0io0l0IoloioOii0oIioOi0[63:0] } ;
 8'h04: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {OL0LLioOOooILOL0LLLIilLl0oLLiIoiL[4*8-1:0] ,O0lIOiilLOiIOollILlioiiOOiiLOO00i[8*8-1:0] ,O0O0oIOiIOLL0LILLIILOOliLO0oO0ilL[8*8-1:0] ,OIiLIoliOIilIl0O00Li00oIO0OlIiooo[31:0] ,OIIli0o0iiLOoOlilIoLIooOIooIL0ilI[63:0] } ;
 8'h08: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {Ol000OloII0LlIII00IIOIlOiioOo0Iii[4*8-1:0] ,OOoOoLoIlLoiILLOlL0ooILOio0OLlI0I[8*8-1:0] ,OOIi0LIIiIoiIIl0OoilO0iIoLloOiIll[8*8-1:0] ,OoOOoIoIoOI0IlllILLlOLOloLoo0IO0I[31:0] ,OllLLOLl0o0Ii0i00lOiLOOOLllIlLoio[63:0] } ;
 8'h10: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {O00I0iOoILll0oILl0ILloii0LIIOOiIO[4*8-1:0] ,OlolloloolOo0o0LLLIl00Li0iiLl00ol[8*8-1:0] ,OIIli0ilooIlOLI0lLO0Oi0IilILOolii[8*8-1:0] ,OlOlIILOLLIll0lo0lO0IOliliOOiL0oI[31:0] ,OoOOLol000OllOLI0LO0LO0LoIliO0iiL[63:0] } ;
 8'h20: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {OO00IIiOlOioiOLIiIloilLII0lLL0OOi[4*8-1:0] ,OOLIlLlLIloIOoooilolooLloIi0OiiIi[8*8-1:0] ,OiiLLiLi0OOlLoOlLOI00ilIL0iLO0lOO[8*8-1:0] ,OiIoI00iOLLOlIiO0I0OlIOL0oLIioIIO[31:0] ,OoLOolIOLlOIIlIiOioiIIOL0lioliOIi[63:0] } ;
 8'h40: OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {OlOl0iOIioolOiill0OLOloOoLiIlllol[4*8-1:0] ,OiIiIlii0O0IIO0oolOlooL0oL0LIIIIO[8*8-1:0] ,OloILiOiLoIOOl0IoloOlI00Oollol0lL[8*8-1:0] ,OiII0LiLIl0OLLIiLIoLlI0l00oLioLoI[31:0] ,OlOIIL0Oi0lLOLl0olL0lLooOIiLioOlI[63:0] } ;
 8'h80 : OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= {OOooOoIiooIliiO0LoLiOlOoIlOOo00I0[4*8-1:0] ,OlIoO0LIi0LOLoLLOoliioiIOolIl00OO[8*8-1:0] ,O0LlLoi0OIilllOOIOl0l0LIOOoLOil0L[8*8-1:0] ,OL0IiIiILoIoIOI0OLOo0l0iOl0OIOlIl[31:0] ,OLLiOOIoo0LlIi0Ll0ol000OIl0LlIiIo[63:0] } ;
 default : OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi <= OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= 256'd0 ;
 OlilIo0olII00llLOlLIloLL0l0iOIOLo <= 1'd0 ;
 end
 else begin
 OlilIo0olII00llLOlLIloLL0l0iOIOLo <= |Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15:8] ;
 case ( Ooli0O0IloLOO0OooL0lIOiiOl000IoO0[15:8]) 8'h01: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {OioOlIooLl0IL0LiioIlILIolO0o0ii0l[4*8-1:0] ,OLllLIi0I0LiLOllOL0ILLlLoLiIOiLoI[8*8-1:0] ,OI0ILilL0olIiOoL0lOiiooolOOllIIIL[8*8-1:0] ,O0000LloLiliiLOoIi0iLiLli0iloOOLI[31:0] ,OOIlLiILIoIiLLLIoIoi0IiIoo0OoIOil[63:0] } ;
 8'h02: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {Ol0i0IoiOlliILloOOlIL0oOOl0LIi0o0[4*8-1:0] ,Oloo0IIooolliliLOLoLoL0oI0LOliLlL[8*8-1:0] ,OIiIIlooOiolooLoI0iLi0loLiloiLOll[8*8-1:0] ,OlLLLIIoliL0Ol0lLLiil0ol0OlolIIIl[31:0] ,OI0IOio0lIIOiLllLLLIoIoiIoiOLillO[63:0] } ;
 8'h04: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {OIIiIl0Oo0OLOoLi0O0Iil0IOO0LiIliO[4*8-1:0] ,O00oIiiOLOoilolOol0OIIOII00lllOIo[8*8-1:0] ,OO0ilOiiOiIooOlIiO0l00iOliILoOIIi[8*8-1:0] ,OoL0IILLIoLlIilIlIoOoiOio0Iol0lLI[31:0] ,Oo0I0llOI0ioOlIio0Io0oIlOlIOlIILI[63:0] } ;
 8'h08: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {OLIIioOL00o0iOlL0l0oLoI0OO0iLoOol[4*8-1:0] ,OlLi0LOI0LoLioI0loilIlo00iliILIoi[8*8-1:0] ,OOiiLOIIOolOIOl0I0LOIlioIIll0iIIO[8*8-1:0] ,OI00ilIioiLo0ioiiIi0O0IolOiOi00IO[31:0] ,OiOoiILoiIiIIoll0loilLl00Ll00O0iL[63:0] } ;
 8'h10: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {OoIIOolLOL0oiOO0O0L0iiLlolIiiOLII[4*8-1:0] ,OLioIOLOILilililoO0ililOi0oiIoo0o[8*8-1:0] ,OLlliOLLil0LiIo0Il0iOOl0lIiIi0loL[8*8-1:0] ,Ool0i0Oliiil000lLLlOiIOLOIOIi0Lll[31:0] ,Oo0IoILIliiOo0oooOLOiIo00i0L00Iio[63:0] } ;
 8'h20: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {OoLO0LoiiIL0lilol0oloO0loiLLiIIl0[4*8-1:0] ,OLI0OlLLOll0LooOOiLIlOLoIoiLOO0oL[8*8-1:0] ,OoOLolo0o0IOilOOLI0OoioLilIliI0lO[8*8-1:0] ,O0o0OiliollLIi0IiLilIiOlLOOOLO00i[31:0] ,OOooiloOoOIIiOiiLlLlLlIOIOIlolIol[63:0] } ;
 8'h40: OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {O0oOL0illOloooo0ioIiOLOooLILllLl0[4*8-1:0] ,Oloo0LO0LL0Io0l00lLLLIolI0lIlLiLo[8*8-1:0] ,OlOL0OLLooilLiOliIOIOOlIio00Oiili[8*8-1:0] ,OO0oolOlI0iloil0ooIolIioiol00I00I[31:0] ,O0oo0ILLOL0ioL0LIOiOiLIL0iol0ooiI[63:0] } ;
 8'h80 : OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= {OLiILioillIololIOILoOLlI0LILLliIL[4*8-1:0] ,OoOOillllIiloIOIILO0lL0LIl0iOlIII[8*8-1:0] ,OoiLiIoIIIiOo0O0OoI0oOi0OOiOOliLi[8*8-1:0] ,OLIoIliI0LI0liL0i0IIIiLloL000l0lO[31:0] ,Oo00OloiOIoLi00Oo0ooiololoOoooLLO[63:0] } ;
 default : OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 <= OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0000Lil0OoOOILlIlOlooioiIOloOioi <= 256'd0 ;
 end
 else if ( OLLliiOoIi0oLoIlllooooiLIoLOlL0iO ) begin
 O0000Lil0OoOOILlIlOlooioiIOloOioi <= OLoI0oOO00OoL0LiIOi0LLOlIIIoLoIoi ;
 end
 else if ( OilL0oiOIollIOIOOO0I0IIoLLOoOOOLO ) begin
 O0000Lil0OoOOILlIlOlooioiIOloOioi <= OiILLiLiIiIlIlIOloOlIoOOollIlOiio ;
 end
 else if ( OlilIo0olII00llLOlLIloLL0l0iOIOLo ) begin
 O0000Lil0OoOOILlIlOlooioiIOloOioi <= OIOolOLllIolOllo0lI0iLIo0O0IiLiL0 ;
 end
 else if ( O0i0oLliiiIoIi0iIi00ILlIooi0OLlil ) begin
 O0000Lil0OoOOILlIlOlooioiIOloOioi <= OooiiLl0L0OoiIoi0lo0iIIlLiLlioLIi ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O00lOOl0oILIoiioLOOI0OoioILioLiiL <= 32'd0 ;
 end
 else begin
 case ({O0i00oOl00OoIIOIil0LLOi0looIOIL00,Ooli0O0IloLOO0OooL0lIOiiOl000IoO0}) 33'h0_0000_0001: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {Ooii00l0ooOoIliILL0lLLLLLoILlIIoO[31:0]} ;
 33'h0_0000_0002: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OILl0LOii0lOi0LlLIIoIL0LLOoli0oll[31:0]} ;
 33'h0_0000_0004: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {O0Io0oIliooLo0i0i0lL0IlILOloiiIlI[31:0]} ;
 33'h0_0000_0008: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OLLli0LLl0LlILOoi000iLoiiOOOLooLI[31:0]} ;
 33'h0_0000_0010: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OoIooi0LILolioIilliiol0I0iLoioIoi[31:0]} ;
 33'h0_0000_0020: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OILolilliOIlLILOoioLii0iI0lII0oil[31:0]} ;
 33'h0_0000_0040: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OOIilioOiLLoOIL0iLoILiLLliiio0LOl[31:0]} ;
 33'h0_0000_0080: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OiIiOI0iOiOLlLooo0i0O0ilOIoloIL0l[31:0]} ;
 33'h0_0000_0100: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OllioLi0iLLoIOlILoIL0oOO0OiIliOOi[31:0]} ;
 33'h0_0000_0200: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OlOoOLLlO0LOilOiiOoiOi0o0lollolLl[31:0]} ;
 33'h0_0000_0400: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OILoioOioIOL0lIOLoIlIOlolLiOLlIoo[31:0]} ;
 33'h0_0000_0800: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OoI0i0iiiL0ililIOLiL0IioLIL0IooOo[31:0]} ;
 33'h0_0000_1000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OioIoIoo0iIIlOilLlIoILioo0I0lo00o[31:0]} ;
 33'h0_0000_2000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OIIOOi0ilOiLO0ooIo00iOoIo0OIl0il0[31:0]} ;
 33'h0_0000_4000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OLI00Il0O0lI0OoLI0oIloiOIiiILIill[31:0]} ;
 33'h0_0000_8000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {Ooii00oOIo0LioI0lLiIiLI0oooOiiLoL[31:0]} ;
 33'h0_0001_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OioOiiiOlioLLOllo0IiIOiOOli0oi0LI[31:0]} ;
 33'h0_0002_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {O0i000LoOoll00lolOOOOIO0Oio0LIO0o[31:0]} ;
 33'h0_0004_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {Oi0Ol0lLIi00LiiLOoIlIIlIoII0OlOiO[31:0]} ;
 33'h0_0008_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OIlOooOloOi0oL0IoIiOo0lilLIIiLOIl[31:0]} ;
 33'h0_0010_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {Oiio0oo000ioIO0llioIoLILlIlIOOloL[31:0]} ;
 33'h0_0020_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OIooL0lILLIloiOOLiI0ilOIli0LOL000[31:0]} ;
 33'h0_0040_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OILlOiiL00II0oiOlOoOI0lI00I0oIIIi[31:0]} ;
 33'h0_0080_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OLoOiiL00iolo0LOliOll0I0ILIOL0iLI[31:0]} ;
 33'h0_0100_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OII0Iill0IOLO000li0iL0iLoiIoOoliL[31:0]} ;
 33'h0_0200_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OOI0I0II0oOOO0LiLoO0I00LloOllilIl[31:0]} ;
 33'h0_0400_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OOIioIlLoOL00lOliIIllL00illo0L00o[31:0]} ;
 33'h0_0800_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OLiloooloollOoil0LlolLolOILlO00Ol[31:0]} ;
 33'h0_1000_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OOilLILioilLIliOlOoilOOIolLLiLl0I[31:0]} ;
 33'h0_2000_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OlO0loIioIiOiLI0LLLLiLOLlOiiOo0I0[31:0]} ;
 33'h0_4000_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OOlLOll0O0OoL0L0oLlIiiOiOL0o0OoOI[31:0]} ;
 33'h0_8000_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {OIiLOlOll0ol0OOLIo0oOiIilII0Io00L[31:0]} ;
 33'h1_0000_0000: O00lOOl0oILIoiioLOOI0OoioILioLiiL <= {O0liLooiLliIoLOllliIlo0ILo0I0oOOl[31:0] } ;
 default : O00lOOl0oILIoiioLOOI0OoioILioLiiL <= O00lOOl0oILIoiioLOOI0OoioILioLiiL ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0iioiILo0ol0ollLilLl0lO0oI0ilOiL <= 1'd0 ;
 end
 else if (O0i00oOl00OoIIOIil0LLOi0looIOIL00|| (|Ooli0O0IloLOO0OooL0lIOiiOl000IoO0) ) begin
 O0iioiILo0ol0ollLilLl0lO0oI0ilOiL <= 1'd1 ;
 end
 else if ( O0iioiILo0ol0ollLilLl0lO0oI0ilOiL &&(OLILoI0O0oiLILloooL0OLL0iOIoiIoIo==2'd3)) begin
 O0iioiILo0ol0ollLilLl0lO0oI0ilOiL <= 1'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLILoI0O0oiLILloooL0OLL0iOIoiIoIo <= 2'd0 ;
 end
 else if ( O0iioiILo0ol0ollLilLl0lO0oI0ilOiL ) begin
 OLILoI0O0oiLILloooL0OLL0iOIoiIoIo <= OLILoI0O0oiLILloooL0OLL0iOIoiIoIo + 1'd1 ;
 end
 else begin
 OLILoI0O0oiLILloooL0OLL0iOIoiIoIo <= 2'd0 ;
 end
 end
 endmodule
 `timescale 1ns/1ns module OoLiL0iillLiLlLlO0loIIoLl0l0l0LoI ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI , OOiiILlloiOoI0OlilIOoiiLOOLol0IoI , OI00OiLolooiIIiiILoIliO0O0loolIlI , O0Loo0iiI0OlLOlOIiILOooOOlIoioOli , O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo , OILIloOoilLIL00IIOoOilLOO0L0iiIOO , O0oLLi0Ill00l0lioiLioiooIllloIiIl , OilOIloOO0LiLoIL0IIILoIi0Loilll0I , Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 , OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O , OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO , OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 , OlOI0loIIIlOi0OOloOioOIo0L00iOiOi , OO0LlIOOoILoolO0LlO0O0liOIl0OiOil , OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL , OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 , OiooiLLioLLL0lII00ol0oIOllLlOiLlL , OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi , O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 , Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO , O0i0IiOL0liOOoLoOiioLOiIIioolOlLI , OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o , OilLIO0lI0LO0LolOOilILl0oiIlolOlo , OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O , OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL , OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 , OlIIIILlOLoIIio0lIloiiLOIOoliL0IO , OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO , OIoliiOo0i000ooilOOLOiil0LlLiOoLo , Oo00OlooOo0io0OoIloiioLiOlL0llio0 , OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL , OOoOoILioOoIlIoLliOLOOi0io0IlLolo , OiLllooo0Li0lioiolLi0ILIoLOliil0I , OlioIL00LLooOiOiOi0liiLI0OOLLI0lO , OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl , OlIlI0o0I0ILOloiOioI0i0IiIliLil00 , OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo , OLL0OiLILloil0IoOlLIIloLIiIlllLil , OILI0LLillilOlllLil0ioLoIiliOoLLo , OiIOlO00OOiiOlOloOOIl0IIoL00IOliL , OoIloII0oLiOLOLIllOL0iOoooOliOIii , Ol0iOoOil0il0LilI0Io0IIooll0i0I0o , OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL , O0oill0llILOilo0i0LIoOLIoolL0Il0o , OlliILlLOilOl0LO0O0OilooiIIiOi0Ll , OiL0LolLLIOlliloII00llOil0oIlOiIo , O0llIOIliLOO0iiOoO0OO0lIOloLoII0I , OOLoL0looIOoioIoOooIoLIiIiLiLoiOl , OIoIooIolOilIOlooOlOIIOoilLioOIIO , Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l , O0IOooLliOlIllOliILoolIIoIiO0Ilol , OolIOLOooiLLIllI0LOLIolllLoilolIl , OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 , O0lOIlooLi0lilOllLlilIo00iOLiOLLo , Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI );
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input [31:0] OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ;
 input [31:0] OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ;
 input [31:0] OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 input O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ;
 output [31:0] OilOIloOO0LiLoIL0IIILoIi0Loilll0I ;
 output [31:0] Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 ;
 output [31:0] OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ;
 output [63:0] OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ;
 output [ 2:0] OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ;
 output [ 2:0] OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ;
 output [ 2:0] OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ;
 output [ 2:0] OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ;
 output [ 2:0] OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ;
 output [ 2:0] OiooiLLioLLL0lII00ol0oIOllLlOiLlL ;
 output [ 2:0] OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ;
 output [ 2:0] O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ;
 output [ 2:0] Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ;
 output [ 2:0] O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ;
 output [ 2:0] OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ;
 output [ 2:0] OilLIO0lI0LO0LolOOilILl0oiIlolOlo ;
 output [ 2:0] OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ;
 output [ 2:0] OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ;
 output [ 2:0] OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ;
 output [ 2:0] OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ;
 output [ 2:0] OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ;
 output [ 2:0] OIoliiOo0i000ooilOOLOiil0LlLiOoLo ;
 output [ 2:0] Oo00OlooOo0io0OoIloiioLiOlL0llio0 ;
 output [ 2:0] OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ;
 output [ 2:0] OOoOoILioOoIlIoLliOLOOi0io0IlLolo ;
 output [ 2:0] OiLllooo0Li0lioiolLi0ILIoLOliil0I ;
 output [ 2:0] OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ;
 output [ 2:0] OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ;
 output [ 2:0] OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ;
 output [ 2:0] OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ;
 output [ 2:0] OLL0OiLILloil0IoOlLIIloLIiIlllLil ;
 output [ 2:0] OILI0LLillilOlllLil0ioLoIiliOoLLo ;
 output [ 2:0] OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ;
 output [ 2:0] OoIloII0oLiOLOLIllOL0iOoooOliOIii ;
 output [ 2:0] Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ;
 output [ 2:0] OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ;
 input O0oill0llILOilo0i0LIoOLIoolL0Il0o ;
 input OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ;
 input OiL0LolLLIOlliloII00llOil0oIlOiIo ;
 input O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ;
 input [ 5:0] Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 input OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ;
 input OIoIooIolOilIOlooOlOIIOoilLioOIIO ;
 input [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 input [ 15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 input OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 input [191:0] O0lOIlooLi0lilOllLlilIo00iOLiOLLo ;
 input [ 15:0] O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ;
 input [ 15:0] OILIloOoilLIL00IIOoOilLOO0L0iiIOO ;
 input [ 31:0] O0oLLi0Ill00l0lioiLioiooIllloIiIl ;
 reg [31:0] OilOIloOO0LiLoIL0IIILoIi0Loilll0I ;
 reg [31:0] OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O ;
 reg [63:0] OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO ;
 reg [ 2:0] OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 ;
 reg [ 2:0] OlOI0loIIIlOi0OOloOioOIo0L00iOiOi ;
 reg [ 2:0] OO0LlIOOoILoolO0LlO0O0liOIl0OiOil ;
 reg [ 2:0] OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL ;
 reg [ 2:0] OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 ;
 reg [ 2:0] OiooiLLioLLL0lII00ol0oIOllLlOiLlL ;
 reg [ 2:0] OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi ;
 reg [ 2:0] O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 ;
 reg [ 2:0] Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO ;
 reg [ 2:0] O0i0IiOL0liOOoLoOiioLOiIIioolOlLI ;
 reg [ 2:0] OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o ;
 reg [ 2:0] OilLIO0lI0LO0LolOOilILl0oiIlolOlo ;
 reg [ 2:0] OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O ;
 reg [ 2:0] OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL ;
 reg [ 2:0] OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 ;
 reg [ 2:0] OlIIIILlOLoIIio0lIloiiLOIOoliL0IO ;
 reg [ 2:0] OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO ;
 reg [ 2:0] OIoliiOo0i000ooilOOLOiil0LlLiOoLo ;
 reg [ 2:0] Oo00OlooOo0io0OoIloiioLiOlL0llio0 ;
 reg [ 2:0] OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL ;
 reg [ 2:0] OOoOoILioOoIlIoLliOLOOi0io0IlLolo ;
 reg [ 2:0] OiLllooo0Li0lioiolLi0ILIoLOliil0I ;
 reg [ 2:0] OlioIL00LLooOiOiOi0liiLI0OOLLI0lO ;
 reg [ 2:0] OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl ;
 reg [ 2:0] OlIlI0o0I0ILOloiOioI0i0IiIliLil00 ;
 reg [ 2:0] OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo ;
 reg [ 2:0] OLL0OiLILloil0IoOlLIIloLIiIlllLil ;
 reg [ 2:0] OILI0LLillilOlllLil0ioLoIiliOoLLo ;
 reg [ 2:0] OiIOlO00OOiiOlOloOOIl0IIoL00IOliL ;
 reg [ 2:0] OoIloII0oLiOLOLIllOL0iOoooOliOIii ;
 reg [ 2:0] Ol0iOoOil0il0LilI0Io0IIooll0i0I0o ;
 reg [ 2:0] OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL ;
 wire [31:0] Ol0oLlOIoOl0iLLLiilOI0ioo0iIoLLo0 = 32'd0 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I <= 32'd0 ;
 end
 else if ( O0oill0llILOilo0i0LIoOLIoolL0Il0o && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 0] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 1] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 2] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 3] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 4] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 5] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 6] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 7] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 8] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 9] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[10] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[11] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[12] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[13] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[14] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[15] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[16] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[17] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[18] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[19] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[20] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[21] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[22] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[23] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[24] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[25] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[26] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[27] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[28] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[29] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[30] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30];
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[31] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31];
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && ( OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4) ) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli && (OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 0] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 1] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 2] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 3] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 4] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 5] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 6] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 7] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 8] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[ 9] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[10] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[11] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[12] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[13] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[14] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[15] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[16] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[17] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[18] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[19] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[20] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[21] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[22] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[23] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[24] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[25] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[26] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[27] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[28] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[29] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[30] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ;
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I[31] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ;
 end
 else begin
 OilOIloOO0LiLoIL0IIILoIi0Loilll0I <= 32'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O <= 32'd0 ;
 end
 else if ( O0oill0llILOilo0i0LIoOLIoolL0Il0o && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 0] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 1] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 2] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 3] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 4] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 5] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 6] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 7] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 8] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 9] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31];
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && ( OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4) ) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 0] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 1] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 2] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 3] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 4] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 5] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 6] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 7] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 8] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 9] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ;
 end
 else if ( OOLoL0looIOoioIoOooIoLIiIiLiLoiOl && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 0] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 1] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 2] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 3] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 4] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 5] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 6] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 7] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 8] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 9] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31];
 end
 else if ( OIoIooIolOilIOlooOlOIIOoilLioOIIO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 0] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 1] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 2] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 3] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 4] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 5] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 6] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 7] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 8] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 9] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30];
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] <= OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31];
 end
 else if ( OiL0LolLLIOlliloII00llOil0oIlOiIo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 0] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 0] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 1] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 1] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 2] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 2] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 3] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 3] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 4] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 4] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 5] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 5] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 6] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 6] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 7] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 7] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 8] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 8] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 9] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 9] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[10] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[11] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[12] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[13] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[14] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[15] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[16] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[17] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[18] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[19] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[20] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[21] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[22] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[23] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[24] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[25] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[26] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[27] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[28] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[29] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[30] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[31] ;
 end
 else if ( O0llIOIliLOO0iiOoO0OO0lIOloLoII0I && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>= Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l[5:0] ) ) begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 0] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 0] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 1] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 1] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 2] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 2] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 3] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 3] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 4] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 4] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 5] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 5] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 6] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 6] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 7] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 7] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 8] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 8] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[ 9] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 9] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[10] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[10] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[11] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[11] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[12] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[12] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[13] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[13] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[14] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[14] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[15] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[15] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[16] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[16] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[17] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[17] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[18] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[18] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[19] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[19] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[20] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[20] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[21] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[21] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[22] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[22] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[23] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[23] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[24] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[24] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[25] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[25] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[26] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[26] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[27] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[27] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[28] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[28] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[29] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[29] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[30] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[30] ;
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O[31] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[31] ;
 end
 else begin
 OllIOIIOiLO0OOLl0I0I0LL0OOl0oll0O <= 32'd0 ;
 end
 end
 wire [63: 0] OlIlIOiiLi0llOL0OIioIOI0lILOolOlI = O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64:64+64];
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO <= 64'd0 ;
 end
 else if ( O0oill0llILOilo0i0LIoOLIoolL0Il0o && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO <= OlIlIOiiLi0llOL0OIioIOI0lILOolOlI ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO <= OlIlIOiiLi0llOL0OIioIOI0lILOolOlI ;
 end
 else if ( ( OOLoL0looIOoioIoOooIoLIiIiLiLoiOl || OiL0LolLLIOlliloII00llOil0oIlOiIo) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO <= OlIlIOiiLi0llOL0OIioIOI0lILOolOlI ;
 end
 else if ( OIoIooIolOilIOlooOlOIIOoilLioOIIO && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO <= OlIlIOiiLi0llOL0OIioIOI0lILOolOlI ;
 end
 else if ( O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ) begin
 OilOLLl0LOOliOoLio0lIiI0OoOLLoIOO <= OlIlIOiiLi0llOL0OIioIOI0lILOolOlI ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 <= 3'd0 ;
 OlOI0loIIIlOi0OOloOioOIo0L00iOiOi <= 3'd0 ;
 OO0LlIOOoILoolO0LlO0O0liOIl0OiOil <= 3'd0 ;
 OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL <= 3'd0 ;
 OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 <= 3'd0 ;
 OiooiLLioLLL0lII00ol0oIOllLlOiLlL <= 3'd0 ;
 OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi <= 3'd0 ;
 O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 <= 3'd0 ;
 Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO <= 3'd0 ;
 O0i0IiOL0liOOoLoOiioLOiIIioolOlLI <= 3'd0 ;
 OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o <= 3'd0 ;
 OilLIO0lI0LO0LolOOilILl0oiIlolOlo <= 3'd0 ;
 OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O <= 3'd0 ;
 OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL <= 3'd0 ;
 OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 <= 3'd0 ;
 OlIIIILlOLoIIio0lIloiiLOIOoliL0IO <= 3'd0 ;
 OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO <= 3'd0 ;
 OIoliiOo0i000ooilOOLOiil0LlLiOoLo <= 3'd0 ;
 Oo00OlooOo0io0OoIloiioLiOlL0llio0 <= 3'd0 ;
 OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL <= 3'd0 ;
 OOoOoILioOoIlIoLliOLOOi0io0IlLolo <= 3'd0 ;
 OiLllooo0Li0lioiolLi0ILIoLOliil0I <= 3'd0 ;
 OlioIL00LLooOiOiOi0liiLI0OOLLI0lO <= 3'd0 ;
 OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl <= 3'd0 ;
 OlIlI0o0I0ILOloiOioI0i0IiIliLil00 <= 3'd0 ;
 OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo <= 3'd0 ;
 OLL0OiLILloil0IoOlLIIloLIiIlllLil <= 3'd0 ;
 OILI0LLillilOlllLil0ioLoIiliOoLLo <= 3'd0 ;
 OiIOlO00OOiiOlOloOOIl0IIoL00IOliL <= 3'd0 ;
 OoIloII0oLiOLOLIllOL0iOoooOliOIii <= 3'd0 ;
 Ol0iOoOil0il0LilI0Io0IIooll0i0I0o <= 3'd0 ;
 OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL <= 3'd0 ;
 end
 else if ( (O0oill0llILOilo0i0LIoOLIoolL0Il0o || OIoIooIolOilIOlooOlOIIOoilLioOIIO) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlOI0loIIIlOi0OOloOioOIo0L00iOiOi <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OO0LlIOOoILoolO0LlO0O0liOIl0OiOil <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OiooiLLioLLL0lII00ol0oIOllLlOiLlL <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 O0i0IiOL0liOOoLoOiioLOiIIioolOlLI <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OilLIO0lI0LO0LolOOilILl0oiIlolOlo <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlIIIILlOLoIIio0lIloiiLOIOoliL0IO <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OIoliiOo0i000ooilOOLOiil0LlLiOoLo <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 Oo00OlooOo0io0OoIloiioLiOlL0llio0 <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OOoOoILioOoIlIoLliOLOOi0io0IlLolo <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OiLllooo0Li0lioiolLi0ILIoLOliil0I <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlioIL00LLooOiOiOi0liiLI0OOLLI0lO <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OlIlI0o0I0ILOloiOioI0i0IiIliLil00 <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OLL0OiLILloil0IoOlLIIloLIiIlllLil <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OILI0LLillilOlllLil0ioLoIiliOoLLo <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OiIOlO00OOiiOlOloOOIl0IIoL00IOliL <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OoIloII0oLiOLOLIllOL0iOoooOliOIii <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 Ol0iOoOil0il0LilI0Io0IIooll0i0I0o <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL <= 4'd8 - OolIOLOooiLLIllI0LOLIolllLoilolIl[3:0] ;
 end
 else begin
 OLL00iLoOL0oLOOOOLOloiiLO00i0Ill0 <= 3'd0 ;
 OlOI0loIIIlOi0OOloOioOIo0L00iOiOi <= 3'd0 ;
 OO0LlIOOoILoolO0LlO0O0liOIl0OiOil <= 3'd0 ;
 OlOIOoO0iIi0oolL0i0LoIoilIiiLl0LL <= 3'd0 ;
 OLI0o0ooOOL0LiLOLOoLIIoLiiIOIOoi0 <= 3'd0 ;
 OiooiLLioLLL0lII00ol0oIOllLlOiLlL <= 3'd0 ;
 OlOIOIo0lLIiIlOiIIlIlIIiiLOlioiOi <= 3'd0 ;
 O0i0OlL0IOLiO0lILO0oo0IlLIIoi0oL0 <= 3'd0 ;
 Ololo0OO0iOLIOi0IilIoiOOiIiIoOlOO <= 3'd0 ;
 O0i0IiOL0liOOoLoOiioLOiIIioolOlLI <= 3'd0 ;
 OIIOo0IiL0liOIilOOIoLiIOLOlILOL0o <= 3'd0 ;
 OilLIO0lI0LO0LolOOilILl0oiIlolOlo <= 3'd0 ;
 OiOLOoLoL0o0iiO0Ol0lOiOIOLi0Ill0O <= 3'd0 ;
 OLOOLlLLOilooiOOILiIO0oiOOI0I0LlL <= 3'd0 ;
 OoOl00LoLOllOoO0Ll0iOoO0L00llOOO0 <= 3'd0 ;
 OlIIIILlOLoIIio0lIloiiLOIOoliL0IO <= 3'd0 ;
 OO0iiLLlIil0lILLoLiL0i0LO00iLoiIO <= 3'd0 ;
 OIoliiOo0i000ooilOOLOiil0LlLiOoLo <= 3'd0 ;
 Oo00OlooOo0io0OoIloiioLiOlL0llio0 <= 3'd0 ;
 OooOO0lLol0OO0OiO0IlLIi0LOOLL0ioL <= 3'd0 ;
 OOoOoILioOoIlIoLliOLOOi0io0IlLolo <= 3'd0 ;
 OiLllooo0Li0lioiolLi0ILIoLOliil0I <= 3'd0 ;
 OlioIL00LLooOiOiOi0liiLI0OOLLI0lO <= 3'd0 ;
 OlIIi0iOoIooOI0o0OOlOOIlo0ILllIIl <= 3'd0 ;
 OlIlI0o0I0ILOloiOioI0i0IiIliLil00 <= 3'd0 ;
 OI0LoliIO0oOo0I0Ooo0loIIIIiO0LiOo <= 3'd0 ;
 OLL0OiLILloil0IoOlLIIloLIiIlllLil <= 3'd0 ;
 OILI0LLillilOlllLil0ioLoIiliOoLLo <= 3'd0 ;
 OiIOlO00OOiiOlOloOOIl0IIoL00IOliL <= 3'd0 ;
 OoIloII0oLiOLOLIllOL0iOoooOliOIii <= 3'd0 ;
 Ol0iOoOil0il0LilI0Io0IIooll0i0I0o <= 3'd0 ;
 OIIOOLlOoI0iL0iOoil0ooLIL0LliiLiL <= 3'd0 ;
 end
 end
 endmodule
 module OLiIILolLli0LiLoOOo0lIlOiOoO0lioL ( OOLIiil0IlIllLollIl0LIilliOI0iolo , OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI , OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII , OOLOoolOi0LIo0olO0loLllIlllIiiIiI , OOOLiLOilooIi0Iio00ilILoLIILOoOoI , OLLOooI0ILL00ILloiliILLLiioooLliI , OL0O0IIio0loL0L0Il0li0i00lliIoOOI , OILoli0OIOIIOI0OiliOo0i0OLoliOOiI , Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII , O0lOIlooLi0lilOllLlilIo00iOLiOLLo , O0IOooLliOlIllOliILoolIIoIiO0Ilol , Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl , O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI , O0il0IO0olIoLiOIL0000lo0OoliIL0Ll , Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI );
 input [4:0] OOLIiil0IlIllLollIl0LIilliOI0iolo ;
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ;
 input [ 3:0] OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 input OOLOoolOi0LIo0olO0loLllIlllIiiIiI ;
 input OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 input [63:0] OLLOooI0ILL00ILloiliILLLiioooLliI ;
 input [2:0] OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 input OL0O0IIio0loL0L0Il0li0i00lliIoOOI ;
 input Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ;
 output [191:0] O0lOIlooLi0lilOllLlilIo00iOLiOLLo ;
 output [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 input [ 5:0] Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ;
 input O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ;
 output O0il0IO0olIoLiOIL0000lo0OoliIL0Ll ;
 reg [191:0] O0lOIlooLi0lilOllLlilIo00iOLiOLLo ;
 reg [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol;
 wire [ 5:0] Oll0iI00Ii0IiiOoo0ioLilOiIL0i0LIO ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0IOooLliOlIllOliILoolIIoIiO0Ilol <= 6'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 O0IOooLliOlIllOliILoolIIoIiO0Ilol <= 6'd8 - OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII - OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 end
 else if (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII) begin
 O0IOooLliOlIllOliILoolIIoIiO0Ilol <= 6'd0 ;
 end
 else if ( (OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI)&&(O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI) ) begin
 O0IOooLliOlIllOliILoolIIoIiO0Ilol <= O0IOooLliOlIllOliILoolIIoIiO0Ilol + 6'd8 - Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl - OILoli0OIOIIOI0OiliOo0i0OLoliOOiI;
 end
 else if ( OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI ) begin
 O0IOooLliOlIllOliILoolIIoIiO0Ilol <= O0IOooLliOlIllOliILoolIIoIiO0Ilol + 6'd8 - OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 end
 else if ( O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ) begin
 O0IOooLliOlIllOliILoolIIoIiO0Ilol <= O0IOooLliOlIllOliILoolIIoIiO0Ilol - Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ;
 end
 end
 assign Oll0iI00Ii0IiiOoo0ioLilOiIL0i0LIO = O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? ( O0IOooLliOlIllOliILoolIIoIiO0Ilol-Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ) : O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 reg [191:0] OioLil0Iili0llOliOIooOiOlO0iii0LI;
 wire [191:0] OillLiOl0Llil0o0OiLo0L0oiLOOiIILO;
 reg [191:0] OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO;
 wire [191:0] Olil0I0oIiLiooIIIILIoiIio0iI0L0Ii;
 assign OillLiOl0Llil0o0OiLo0L0oiLOOiIILO = O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? OioLil0Iili0llOliOIooOiOlO0iii0LI : O0lOIlooLi0lilOllLlilIo00iOLiOLLo ;
 always@ (*) begin
 case ( Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ) 5'd0 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[127+64: 0] } ;
 5'd1 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[119+64: 0] , 8'd0 } ;
 5'd2 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[111+64: 0] , 16'd0 } ;
 5'd3 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[103+64: 0] , 24'd0 } ;
 5'd4 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 95+64: 0] , 32'd0 } ;
 5'd5 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 87+64: 0] , 40'd0 } ;
 5'd6 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 79+64: 0] , 48'd0 } ;
 5'd7 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 71+64: 0] , 56'd0 } ;
 5'd8 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63+64: 0] , 64'd0 } ;
 5'd9 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 55+64: 0] , 72'd0 } ;
 5'd10 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 47+64: 0] , 80'd0 } ;
 5'd11 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 39+64: 0] , 88'd0 } ;
 5'd12 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 31+64: 0] , 96'd0 } ;
 5'd13 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 23+64: 0] ,104'd0 } ;
 5'd14 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 15+64: 0] ,112'd0 } ;
 5'd15 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 7+64: 0] ,120'd0 } ;
 5'd16 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 63: 0] ,128'd0 } ;
 5'd17 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 55: 0] ,136'd0 } ;
 5'd18 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 47: 0] ,144'd0 } ;
 5'd19 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 39: 0] ,152'd0 } ;
 5'd20 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 31: 0] ,160'd0 } ;
 5'd21 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 23: 0] ,168'd0 } ;
 5'd22 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 15: 0] ,176'd0 } ;
 5'd23 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { O0lOIlooLi0lilOllLlilIo00iOLiOLLo[ 7: 0] ,184'd0 } ;
 5'd24 : OioLil0Iili0llOliOIooOiOlO0iii0LI = { 192'd0 } ;
 default : OioLil0Iili0llOliOIooOiOlO0iii0LI = { 192'd0 } ;
 endcase end
 always@ (*) begin
 case ( Oll0iI00Ii0IiiOoo0ioLilOiIL0i0LIO ) 5'd0 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] ,128'd0 } ;
 5'd1 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64:120+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] ,120'd0 } ;
 5'd2 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64:112+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] ,112'd0 } ;
 5'd3 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64:104+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] ,104'd0 } ;
 5'd4 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 96+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 96'd0 } ;
 5'd5 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 88+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 88'd0 } ;
 5'd6 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 80+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 80'd0 } ;
 5'd7 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 72+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 72'd0 } ;
 5'd8 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 64+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 64'd0 } ;
 5'd9 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 56+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 56'd0 } ;
 5'd10 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 48+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 48'd0 } ;
 5'd11 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 40+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 40'd0 } ;
 5'd12 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 32+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 32'd0 } ;
 5'd13 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 24+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 24'd0 } ;
 5'd14 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 16+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 16'd0 } ;
 5'd15 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 8+64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] , 8'd0 } ;
 5'd16 : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] } ;
 default : OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO = { OillLiOl0Llil0o0OiLo0L0oiLOOiIILO[127+64: 64],OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] } ;
 endcase end
 assign Olil0I0oIiLiooIIIILIoiIio0iI0L0Ii = OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI ? OOLoIOllILIOo0iOiLOOo0I0oLL0ioiiO : OillLiOl0Llil0o0OiLo0L0oiLOOiIILO ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= 192'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 case ( OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ) 3'd0 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[63:0] ,64'd0 ,64'd0 } ;
 3'd1 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[55:0] , 8'd0 ,64'd0 ,64'd0 } ;
 3'd2 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[47:0] , 16'd0 ,64'd0 ,64'd0 } ;
 3'd3 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[39:0] , 24'd0 ,64'd0 ,64'd0 } ;
 3'd4 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[31:0] , 32'd0 ,64'd0 ,64'd0 } ;
 3'd5 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[23:0] , 40'd0 ,64'd0 ,64'd0 } ;
 3'd6 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[15:0] , 48'd0 ,64'd0 ,64'd0 } ;
 3'd7 : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { OLLOooI0ILL00ILloiliILLLiioooLliI[ 7:0] , 56'd0 ,64'd0 ,64'd0 } ;
 default : O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= { 64'd0 ,64'd0 ,64'd0 } ;
 endcase end
 else if (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII) begin
 O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= 192'd0 ;
 end
 else if ( (OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI) || (O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI) ) begin
 O0lOIlooLi0lilOllLlilIo00iOLiOLLo <= Olil0I0oIiLiooIIIILIoiIio0iI0L0Ii ;
 end
 end
 /* reg [23:0] OOOIiOlOIl0olilOIIIOOlOl0l0LOollO ;
 reg [23:0] OIiIL0LOiIiIILollOLLiioLLolol0oL0 ;
 reg [23:0] OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0;
 wire [23:0] O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO;
 reg [23:0] O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl;
 wire [23:0] OloliiILlOiOiILlli0IOIoio00iO0ioO;
 assign O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO = O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO ;
 always@ (*) begin
 case ( Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ) 6'd0 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 15+8: 0] } ;
 6'd1 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 14+8: 0] , 1'd0 } ;
 6'd2 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 13+8: 0] , 2'd0 } ;
 6'd3 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 12+8: 0] , 3'd0 } ;
 6'd4 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 11+8: 0] , 4'd0 } ;
 6'd5 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 10+8: 0] , 5'd0 } ;
 6'd6 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 9+8: 0] , 6'd0 } ;
 6'd7 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 8+8: 0] , 7'd0 } ;
 6'd8 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 7+8: 0] , 8'd0 } ;
 6'd9 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 6+8: 0] , 9'd0 } ;
 6'd10 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 5+8: 0] ,10'd0 } ;
 6'd11 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 4+8: 0] ,11'd0 } ;
 6'd12 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 3+8: 0] ,12'd0 } ;
 6'd13 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 2+8: 0] ,13'd0 } ;
 6'd14 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 1+8: 0] ,14'd0 } ;
 6'd15 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 8: 0] ,15'd0 } ;
 6'd16 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 7: 0] ,16'd0 } ;
 6'd17 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 6: 0] ,17'd0 } ;
 6'd18 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 5: 0] ,18'd0 } ;
 6'd19 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 4: 0] ,19'd0 } ;
 6'd20 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 3: 0] ,20'd0 } ;
 6'd21 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 2: 0] ,21'd0 } ;
 6'd22 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 1: 0] ,22'd0 } ;
 6'd23 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { OOOIiOlOIl0olilOIIIOOlOl0l0LOollO[ 0] ,23'd0 } ;
 6'd24 : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { 23'd0 } ;
 default : OII0OoLLlll0oL00ooOlO00Ioo0lLOLi0 = { 23'd0 } ;
 endcase end
 always@ (*) begin
 case ( Oll0iI00Ii0IiiOoo0ioLilOiIL0i0LIO ) 5'd0 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { {8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 8'd0 ,8'd0 } ;
 5'd1 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8 ],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 7'd0 ,8'd0 } ;
 5'd2 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8:14+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 6'd0 ,8'd0 } ;
 5'd3 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8:13+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 5'd0 ,8'd0 } ;
 5'd4 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8:12+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 4'd0 ,8'd0 } ;
 5'd5 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8:11+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 3'd0 ,8'd0 } ;
 5'd6 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8:10+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 2'd0 ,8'd0 } ;
 5'd7 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 9+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} , 1'd0 ,8'd0 } ;
 5'd8 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 8+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,8'd0 } ;
 5'd9 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 7+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,7'd0 } ;
 5'd10 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 6+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,6'd0 } ;
 5'd11 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 5+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,5'd0 } ;
 5'd12 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 4+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,4'd0 } ;
 5'd13 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 3+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,3'd0 } ;
 5'd14 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 2+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,2'd0 } ;
 5'd15 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 1+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} ,1'd0 } ;
 5'd16 : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} } ;
 default : O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl = { O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO[15+8: 8+8],{8{OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI}} } ;
 endcase end
 assign OloliiILlOiOiILlli0IOIoio00iO0ioO = OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI ? O0OLl0iL0oOLOoLiiIiiIOOLL0iL00OLl : O0LiIlollliiOo0IIoIIoIlO0LLo0ooiO ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= 16'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 case ( OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ) 3'd0 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 8'hff , 8'd0,8'd0 } ;
 3'd1 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 7'h7f , 9'd0,8'd0 } ;
 3'd2 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 6'h3f , 10'd0,8'd0 } ;
 3'd3 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 5'h1f , 11'd0,8'd0 } ;
 3'd4 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 4'hf , 12'd0,8'd0 } ;
 3'd5 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 3'h3 , 13'd0,8'd0 } ;
 3'd6 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 2'h2 , 14'd0,8'd0 } ;
 3'd7 : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 1'h1 , 15'd0,8'd0 } ;
 default : OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= { 16'd0,8'd0 } ;
 endcase end
 else if (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII) begin
 OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= 'd0 ;
 end
 else if ( (OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI) || (O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI) ) begin
 OOOIiOlOIl0olilOIIIOOlOl0l0LOollO <= OloliiILlOiOiILlli0IOIoio00iO0ioO ;
 end
 end
 reg [23:0] OiIoolI0Il0i0OILil00iiLllIioolI0O;
 wire [23:0] OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL;
 reg [23:0] OIOliiloIillOoiiooolOoOilLo0oIIoL;
 wire [23:0] OOlolo0OOoLiLl0OiOiooiIOliLlii0lO;
 assign OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL = O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ? OiIoolI0Il0i0OILil00iiLllIioolI0O : OIiIL0LOiIiIILollOLLiioLLolol0oL0 ;
 always@ (*) begin
 case ( Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ) 5'd0 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 15+8: 0] } ;
 5'd1 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 14+8: 0] , 1'd0 } ;
 5'd2 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 13+8: 0] , 2'd0 } ;
 5'd3 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 12+8: 0] , 3'd0 } ;
 5'd4 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 11+8: 0] , 4'd0 } ;
 5'd5 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 10+8: 0] , 5'd0 } ;
 5'd6 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 9+8: 0] , 6'd0 } ;
 5'd7 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 8+8: 0] , 7'd0 } ;
 5'd8 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 7+8: 0] , 8'd0 } ;
 5'd9 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 6+8: 0] , 9'd0 } ;
 5'd10 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 5+8: 0] ,10'd0 } ;
 5'd11 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 4+8: 0] ,11'd0 } ;
 5'd12 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 3+8: 0] ,12'd0 } ;
 5'd13 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 2+8: 0] ,13'd0 } ;
 5'd14 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 1+8: 0] ,14'd0 } ;
 5'd15 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 0+8: 0] ,15'd0 } ;
 5'd16 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 7: 0] ,16'd0 } ;
 6'd17 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 6: 0] ,17'd0 } ;
 6'd18 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 5: 0] ,18'd0 } ;
 6'd19 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 4: 0] ,19'd0 } ;
 6'd20 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 3: 0] ,20'd0 } ;
 6'd21 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 2: 0] ,21'd0 } ;
 6'd22 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 1: 0] ,22'd0 } ;
 6'd23 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { OIiIL0LOiIiIILollOLLiioLLolol0oL0[ 0] ,23'd0 } ;
 6'd24 : OiIoolI0Il0i0OILil00iiLllIioolI0O = { 23'd0 } ;
 default : OiIoolI0Il0i0OILil00iiLllIioolI0O = { 23'd0 } ;
 endcase end
 always@ (*) begin
 case ( Oll0iI00Ii0IiiOoo0ioLilOiIL0i0LIO ) 5'd0 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { {8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 8'd0 ,8'd0 } ;
 5'd1 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8 ],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 7'd0 ,8'd0 } ;
 5'd2 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8:14+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 6'd0 ,8'd0 } ;
 5'd3 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8:13+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 5'd0 ,8'd0 } ;
 5'd4 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8:12+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 4'd0 ,8'd0 } ;
 5'd5 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8:11+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 3'd0 ,8'd0 } ;
 5'd6 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8:10+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 2'd0 ,8'd0 } ;
 5'd7 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 9+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} , 1'd0 ,8'd0 } ;
 5'd8 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 8+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,8'd0 } ;
 5'd9 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 7+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,7'd0 } ;
 5'd10 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 6+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,6'd0 } ;
 5'd11 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 5+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,5'd0 } ;
 5'd12 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 4+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,4'd0 } ;
 5'd13 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 3+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,3'd0 } ;
 5'd14 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 2+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,2'd0 } ;
 5'd15 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 1+8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} ,1'd0 } ;
 5'd16 : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} } ;
 default : OIOliiloIillOoiiooolOoOilLo0oIIoL = { OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL[15+8: 8],{8{OOLOoolOi0LIo0olO0loLllIlllIiiIiI}} } ;
 endcase end
 assign OOlolo0OOoLiLl0OiOiooiIOliLlii0lO = OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI ? OIOliiloIillOoiiooolOoOilLo0oIIoL : OlLliLIiiIi0OiOO0IlOIOOIIILlLILIL ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIiIL0LOiIiIILollOLLiioLLolol0oL0 <= 24'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 OIiIL0LOiIiIILollOLLiioLLolol0oL0 <= {8'h00,8'h00,8'h00} ;
 end
 else if (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII) begin
 OIiIL0LOiIiIILollOLLiioLLolol0oL0 <= 'd0 ;
 end
 else if ( (OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&OL0O0IIio0loL0L0Il0li0i00lliIoOOI) || (O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI) ) begin
 OIiIL0LOiIiIILollOLLiioLLolol0oL0 <= OOlolo0OOoLiLl0OiOiooiIOliLlii0lO ;
 end
 end
 */ reg O0il0IO0olIoLiOIL0000lo0OoliIL0Ll ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0il0IO0olIoLiOIL0000lo0OoliIL0Ll <= 1'd0 ;
 end
 else if (O0IOooLliOlIllOliILoolIIoIiO0Ilol>6'd24) begin
 /* synthesis translate_off */ $display("%m Error buffer is full !!!!! cnt is %d OOLIiil0IlIllLollIl0LIilliOI0iolo is %h \n ", O0IOooLliOlIllOliILoolIIoIiO0Ilol, OOLIiil0IlIllLollIl0LIilliOI0iolo );
 /* synthesis translate_on */ O0il0IO0olIoLiOIL0000lo0OoliIL0Ll <= 1'd1 ;
 end
 else begin
 O0il0IO0olIoLiOIL0000lo0OoliIL0Ll <= 1'd0 ;
 end
 end
 /* synthesis translate_off */ reg [15:0] OlIO000lOoill0Oloi0Oil0IlIOOIiOOL ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OlIO000lOoill0Oloi0Oil0IlIOOIiOOL <= 16'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 OlIO000lOoill0Oloi0Oil0IlIOOIiOOL <= 16'd8 - OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 end
 else if ( OOOLiLOilooIi0Iio00ilILoLIILOoOoI && OL0O0IIio0loL0L0Il0li0i00lliIoOOI ) begin
 OlIO000lOoill0Oloi0Oil0IlIOOIiOOL <= OlIO000lOoill0Oloi0Oil0IlIOOIiOOL + 16'd8 - OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 end
 end
 reg [15:0] OIlOOlI00O00oOIiI0illLI00liILllio ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OIlOOlI00O00oOIiI0illLI00liILllio <= 16'd0 ;
 end
 else if (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI) begin
 OIlOOlI00O00oOIiI0illLI00liILllio <= 16'd0 ;
 end
 else if ( O0lioLooO0LoLlOilIiOlLlIiiLlOoLLI ) begin
 OIlOOlI00O00oOIiI0illLI00liILllio <= OIlOOlI00O00oOIiI0illLI00liILllio + Oo0oiiLoolIIILo0OII0LoLI0ILILoLLl ;
 end
 end
 /* synthesis translate_on */ endmodule
 module OLIi0oO0OOIIOllOoo000loIOil0OLi0O ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI , OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL , Oo0OiL0Lll000LlioLiooLOLloiLiliii , OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI , OioiIooIlil0liIiOIi0lLLIllOioioli , OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 , OlLloLOlOi0iIiLIlOlLio000LLOLILli , OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 , OOlILOLoilIOloioiIoOLI0L0ooLO0Lll , OolOlIOiIIoII0ll0IllLoOiIllIilOoO , OOIiiol0IOILiLloOLiLOIIlIIolooOIO , OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO , OILili00ILILlO0LIoLlll0oliLio0liL , OoILoooiioLLiIIIoiIoiOIO0OllIlIlL , OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO , OIiiiIlLolLIoIioOoOolloi0L0loLoIL , OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO , O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II , OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO , OOlO0o0i0Io0IOllLoIloiioiliOOlIII , OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I , O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 , OlOlLO00i0Oiooo0lLollo0IILIlLO0OI , OLLliI0IiOiollllIOOLL0oL0IlllO0oI , OLO00iLliol0LLIOOIIO0IiLIllO0IL0O , O0OII0Ili0ilol00OLOLoiOl0OlLo0liO , OOL0lolilI0oIloIoIIILooo0lOLOlolI , OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll , OIO00IOolLoOoOL0ILI00i0olI0IiiOOo , OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO , OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 , OIoiIlOo00oL0iL0o0iooollLlilLoIIo , Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII , O0oill0llILOilo0i0LIoOLIoolL0Il0o , OlliILlLOilOl0LO0O0OilooiIIiOi0Ll , OOLoL0looIOoioIoOooIoLIiIiLiLoiOl , OIoIooIolOilIOlooOlOIIOoilLioOIIO , OiL0LolLLIOlliloII00llOil0oIlOiIo , O0llIOIliLOO0iiOoO0OO0lIOloLoII0I , OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL , OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo , OolIOLOooiLLIllI0LOLIolllLoilolIl , O0IOooLliOlIllOliILoolIIoIiO0Ilol , O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo , OILIloOoilLIL00IIOoOilLOO0L0iiIOO , O0oLLi0Ill00l0lioiLioiooIllloIiIl , OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 , O0Loo0iiI0OlLOlOIiILOooOOlIoioOli , OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI , OOiiILlloiOoI0OlilIOoiiLOOLol0IoI , Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l , OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI , OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII , OOLOoolOi0LIo0olO0loLllIlllIiiIiI , OOOLiLOilooIi0Iio00ilILoLIILOoOoI , OLLOooI0ILL00ILloiliILLLiioooLliI , OILoli0OIOIIOI0OiliOo0i0OLoliOOiI , O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI , OilOOioILlOIIOL0iioIOIi0oloooOoLl, OI00OiLolooiIIiiILoIliO0O0loolIlI , OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo , OoI0IoiILOOLILioiioIOoOLioiiOlIio , OIIOLLOIlOlLoi0oiOioLilOiioiiliLO , O0OlOIIOOIOIioo00liool0iIiI0I0Lll , O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii , OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l , OIiOIl0O0OLllloOl0oOoLoIllIL0illO , Oi0loi0OllIlIoI0ILloIllILIO0IIo0I , OoLOIol0OLIIiloO0oLoiliOl0LilIolI , OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i , OOloOOOOiILOioIlIOO0oILilOLLL00OO, OOIlIOO0IL0OoLli0IoliIioOOlIILlii , OioOlll0OooLLL0IIIIIli0ollooo0L0L , OooOLOOliIlIOlio00OO0oloLoOi0lliO , OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O , OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI , O0I0oI0I000LllOOI0L0lOlIl000LIioO , OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO , OLlOiiLlLoolliOiO0i0lOloio0L0oL00 , OilOI0i0lloo0Lll000I0OIoIOI0lioiO , OlooiiLooL0L00oIIiioLloiIolOoOlLo , OLo0LOlILllLILOIiiiL0LIlLIoLlO0II , OiiOioOIO00LOOLilooiooo0olO0illo0 , OLl0LoLoii00oiOOoilollii000iIOlOI , OLlil0000Oiil0IOOLiloIlliOoLLol0L , OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI , OO0OOILiO000LOILL0OllLi0l0oliLOo0 , OLiLllIIIlo0llILiLloLOoooOLOilI0l , Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl , OiL0IiiliiioOOLliLiiLILlIOloOLL0L , OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi , OllLOLiIilI0oili000OiLilLioIOoIl0 , OOooI0loOL0iiOIoOili0OOOLLiiIiLOl , OLIIiIIIOILl0loi0lO0IiOoolLIloi00 , OoOillIILLoLoOioLloli0OLILlIOOoLo , OlOlO00LLloOiOolOiOLOIiloLil0L0LI , OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO , OlOLIILoL0ll0oooOo0OIoLoOoiLIolol , OIlLOILiLLo0ol0OLlI0IILilILLLlILO , O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i , Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL , OOiIlillllLOI0oOOoILlol0ILoIoOLil , OOIiO0olO0OLlo0liIoiOioiIO00oOIiL , O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 , OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l , OlolLlliLo0O0l0lOOolL0ioI0O0Li00l , Oo0oI0oLOLlloloiiLIIol0LilOlOIliI , OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo , OoiLlL0oiiIloLOoloIL0oLii00IIIoII , Oo0LLillol0loLIo0iOl0oOLlIOlILoIO , OO0liOO0iOOIioool0OoLliiiI0l0ilOo , OiIOLi00lOILlOOL0oLLloL0io0LoIoOL );
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 input [15:0] OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI ;
 input [15:0] OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL ;
 input [15:0] Oo0OiL0Lll000LlioLiooLOLloiLiliii ;
 input [15:0] OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI ;
 input [15:0] OioiIooIlil0liIiOIi0lLLIllOioioli ;
 input [15:0] OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 ;
 input [15:0] OlLloLOlOi0iIiLIlOlLio000LLOLILli ;
 input [15:0] OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 ;
 input [15:0] OOlILOLoilIOloioiIoOLI0L0ooLO0Lll ;
 input [15:0] OolOlIOiIIoII0ll0IllLoOiIllIilOoO ;
 input [15:0] OOIiiol0IOILiLloOLiLOIIlIIolooOIO ;
 input [15:0] OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO ;
 input [15:0] OILili00ILILlO0LIoLlll0oliLio0liL ;
 input [15:0] OoILoooiioLLiIIIoiIoiOIO0OllIlIlL ;
 input [15:0] OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO ;
 input [15:0] OIiiiIlLolLIoIioOoOolloi0L0loLoIL ;
 input [15:0] OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO ;
 input [15:0] O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II ;
 input [15:0] OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO ;
 input [15:0] OOlO0o0i0Io0IOllLoIloiioiliOOlIII ;
 input [15:0] OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I ;
 input [15:0] O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 ;
 input [15:0] OlOlLO00i0Oiooo0lLollo0IILIlLO0OI ;
 input [15:0] OLLliI0IiOiollllIOOLL0oL0IlllO0oI ;
 input [15:0] OLO00iLliol0LLIOOIIO0IiLIllO0IL0O ;
 input [15:0] O0OII0Ili0ilol00OLOLoiOl0OlLo0liO ;
 input [15:0] OOL0lolilI0oIloIoIIILooo0lOLOlolI ;
 input [15:0] OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll ;
 input [15:0] OIO00IOolLoOoOL0ILI00i0olI0IiiOOo ;
 input [15:0] OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO ;
 input [15:0] OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 ;
 input [15:0] OIoiIlOo00oL0iL0o0iooollLlilLoIIo ;
 input Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII ;
 input O0oill0llILOilo0i0LIoOLIoolL0Il0o ;
 input OlliILlLOilOl0LO0O0OilooiIIiOi0Ll ;
 input OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ;
 input OIoIooIolOilIOlooOlOIIOoilLioOIIO ;
 input OiL0LolLLIOlliloII00llOil0oIlOiIo ;
 input O0llIOIliLOO0iiOoO0OO0lIOloLoII0I ;
 input OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL ;
 input [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 input [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 input [15:0] O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo ;
 input [ 15:0] OILIloOoilLIL00IIOoOilLOO0L0iiIOO ;
 input [ 31:0] O0oLLi0Ill00l0lioiLioiooIllloIiIl ;
 input OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 ;
 input O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ;
 output [31:0] OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ;
 output [15:0] Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 output [31:0] OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ;
 input OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ;
 input [ 3:0] OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 input OOLOoolOi0LIo0olO0loLllIlllIiiIiI ;
 input OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 input [63:0] OLLOooI0ILL00ILloiliILLLiioooLliI ;
 input [ 2:0] OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 input [15:0] O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ;
 input [15:0] OilOOioILlOIIOL0iioIOIi0oloooOoLl;
 input [31:0] OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 input [31:0] OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ;
 output OoI0IoiILOOLILioiioIOoOLioiiOlIio ;
 input [15:0] OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ;
 output O0OlOIIOOIOIioo00liool0iIiI0I0Lll ;
 output [ 3:0] O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii ;
 output OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l ;
 output OIiOIl0O0OLllloOl0oOoLoIllIL0illO ;
 output [63:0] Oi0loi0OllIlIoI0ILloIllILIO0IIo0I ;
 output [ 2:0] OoLOIol0OLIIiloO0oLoiliOl0LilIolI ;
 output [15:0] OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i ;
 output [15:0] OOloOOOOiILOioIlIOO0oILilOLLL00OO;
 output [31:0] OOIlIOO0IL0OoLli0IoliIioOOlIILlii ;
 output OioOlll0OooLLL0IIIIIli0ollooo0L0L ;
 output [15:0] OooOLOOliIlIOlio00OO0oloLoOi0lliO ;
 output [31:0] OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ;
 input [31:0] OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ;
 output [31:0] O0I0oI0I000LllOOI0L0lOlIl000LIioO ;
 input [31:0] OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO ;
 input [31:0] OLlOiiLlLoolliOiO0i0lOloio0L0oL00 ;
 input [31:0] OilOI0i0lloo0Lll000I0OIoIOI0lioiO ;
 input [31:0] OlooiiLooL0L00oIIiioLloiIolOoOlLo ;
 input [31:0] OLo0LOlILllLILOIiiiL0LIlLIoLlO0II ;
 input [31:0] OiiOioOIO00LOOLilooiooo0olO0illo0 ;
 input [31:0] OLl0LoLoii00oiOOoilollii000iIOlOI ;
 input [31:0] OLlil0000Oiil0IOOLiloIlliOoLLol0L ;
 input [31:0] OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI ;
 input [31:0] OO0OOILiO000LOILL0OllLi0l0oliLOo0 ;
 input [31:0] OLiLllIIIlo0llILiLloLOoooOLOilI0l ;
 input [31:0] Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl ;
 input [31:0] OiL0IiiliiioOOLliLiiLILlIOloOLL0L ;
 input [31:0] OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi ;
 input [31:0] OllLOLiIilI0oili000OiLilLioIOoIl0 ;
 input [31:0] OOooI0loOL0iiOIoOili0OOOLLiiIiLOl ;
 input [31:0] OLIIiIIIOILl0loi0lO0IiOoolLIloi00 ;
 input [31:0] OoOillIILLoLoOioLloli0OLILlIOOoLo ;
 input [31:0] OlOlO00LLloOiOolOiOLOIiloLil0L0LI ;
 input [31:0] OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO ;
 input [31:0] OlOLIILoL0ll0oooOo0OIoLoOoiLIolol ;
 input [31:0] OIlLOILiLLo0ol0OLlI0IILilILLLlILO ;
 input [31:0] O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i ;
 input [31:0] Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL ;
 input [31:0] OOiIlillllLOI0oOOoILlol0ILoIoOLil ;
 input [31:0] OOIiO0olO0OLlo0liIoiOioiIO00oOIiL ;
 input [31:0] O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0 ;
 input [31:0] OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l ;
 input [31:0] OlolLlliLo0O0l0lOOolL0ioI0O0Li00l ;
 input [31:0] Oo0oI0oLOLlloloiiLIIol0LilOlOIliI ;
 input [31:0] OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo ;
 input [31:0] OoiLlL0oiiIloLOoloIL0oLii00IIIoII ;
 input [31:0] Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ;
 input [31:0] OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 input OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 output [15:0] OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ;
 reg O0OlOIIOOIOIioo00liool0iIiI0I0Lll ;
 reg [ 3:0] O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii ;
 reg OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l ;
 reg OIiOIl0O0OLllloOl0oOoLoIllIL0illO ;
 reg [63:0] Oi0loi0OllIlIoI0ILloIllILIO0IIo0I ;
 reg [ 2:0] OoLOIol0OLIIiloO0oLoiliOl0LilIolI ;
 reg [15:0] OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i ;
 reg [15:0] OOloOOOOiILOioIlIOO0oILilOLLL00OO;
 reg [31:0] OOIlIOO0IL0OoLli0IoliIioOOlIILlii ;
 reg OioOlll0OooLLL0IIIIIli0ollooo0L0L ;
 reg [15:0] OooOLOOliIlIOlio00OO0oloLoOi0lliO ;
 reg OoI0IoiILOOLILioiioIOoOLioiiOlIio ;
 reg [31:0] OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI ;
 reg [31:0] OioL00ILO0li0IO0LIlIO00lL0I0OllIO ;
 reg [31:0] O0I0oI0I000LllOOI0L0lOlIl000LIioO ;
 reg [31:0] OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ;
 reg [31:0] OLOoliOOlOIIIioiilio0liLil0o0I000 ;
 reg [15:0] OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi ;
 reg [15:0] O0IILIl0LlliiloOOlliilOilioILILOO ;
 reg [15:0] OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI ;
 reg [15:0] OlOO0oILoLOLLLLLllOILOLIilOOLL0oL ;
 reg [15:0] O0oIIIlIIiOILloLo0lLlILLOL0LIO00O ;
 reg [15:0] OLLLiliLlOlI00OOlLoLOL00OLoooLIli ;
 reg [15:0] Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo ;
 reg [15:0] OIlilLLloioioO00IlooIl0IoOoiOOl0o ;
 reg [15:0] OLI0O0LOoiLIooi00li0OllLIilLiOiO0 ;
 reg [15:0] OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO ;
 reg [15:0] OilloOilLL0Loolo00OIlloliiIoIlOLL ;
 reg [15:0] O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 ;
 reg [15:0] O0LoILolI0o00OOoiilOlI0io0O0iiiOi ;
 reg [15:0] OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol ;
 reg [15:0] OLlLi0Olo0oloLLoolIi0IIIOlII0LOll ;
 reg [15:0] OL0OIIiI0loIllilLiIlI0oioI0OloIoL ;
 reg [15:0] OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil ;
 reg [15:0] OOI0I0oiooIoOILIL0oLLL0i0iooOL000 ;
 reg [15:0] O0LL0OoiOLiiII0LooolOliI00oIlIlio ;
 reg [15:0] O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl ;
 reg [15:0] OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO ;
 reg [15:0] OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi ;
 reg [15:0] OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo ;
 reg [15:0] OiLOoilOloiOoo0OloLL0llLOIOoLII0O ;
 reg [15:0] OO0loILiiLolIliIOl0oiloLoioiOLloO ;
 reg [15:0] OIL0iiOloLOLO0IooOilOiooOilOoLilO ;
 reg [15:0] OlolILO0OLo0Oi0LiILii00LOlloiLOi0 ;
 reg [15:0] OL0IoII0L0LLo0IOlLILloi0oi0ilIllI ;
 reg [15:0] O00OiLOI0i0oL0lOOI0liiol0iLIlOlii ;
 reg [15:0] O0IoOI0000OlIo0OoiLll0lilIoOLL0ll ;
 reg [15:0] O0LlIILiOiOioLLoi00lIOi0OI00lOO0I ;
 reg [15:0] O0LOIioI0oLioOILLLOi0I0IO0ILoioLO ;
 reg [15:0] OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo ;
 reg [31:0] OliiILooLoLLIi0IliLO0OO0OOiololoL ;
 reg [31:0] Oll0lolIi00IiOOiIl00OI0OLoIioOLOl ;
 reg [31:0] OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I ;
 reg [31:0] OOOiOlOLli0LLiOOLILIllil0OiLLli0L ;
 reg [31:0] O0LiLoL0IooiOILoioILLLLli00o0LI0I ;
 reg [31:0] OIolIiLOiOLoO00oiliiollllO0l0OloO ;
 reg [31:0] Oil0OiILooLiiioloiiI0oLLlOlLllo0i ;
 reg [31:0] OI0LoL000LIII0lI0LL0LoilIiIlLLiOl ;
 reg [31:0] OoiLi0oolILIllloliLiL0LolIliiLOlo ;
 reg [31:0] OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO ;
 reg [31:0] OioooOOI00ollOl0LiLIl0LIliO00OOii ;
 reg [31:0] OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl ;
 reg [31:0] OoolIOILLooLiOLlLiIoO00OooLLL0LLO ;
 reg [31:0] OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0 ;
 reg [31:0] OoIIliiLlI0OilooiiILLLOL0oII0ILio ;
 reg [31:0] OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i ;
 reg [31:0] OliilLooOIL0lio0OOioLLoLoLOlioIio ;
 reg [31:0] OolioiLoIlIlolO0ooiO0OLOoIlIllIi0 ;
 reg [31:0] OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo ;
 reg [31:0] OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo ;
 reg [31:0] O0iiOolLIl0iOLOiLOOLII00IloOo0li0 ;
 reg [31:0] OLilOOlILoL0oioOOOlOLlOl0li0lIli0 ;
 reg [31:0] OlIIiOliliiioo0LO0I0IIOIiLLooI0lI ;
 reg [31:0] OiOllilOOiI0II0IIilo0IllOOIIIoLii ;
 reg [31:0] OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI ;
 reg [31:0] OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l ;
 reg [31:0] OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0 ;
 reg [31:0] OloOLL0I00I0oIIILLo0Ol0Il0lIILL00 ;
 reg [31:0] OioiIOLioLOlOoliOlLli0i0IolIlOLiL ;
 reg [31:0] OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI ;
 reg [31:0] OiIooILlOili0io0LiiiILIloOi0lIIOl ;
 reg [31:0] OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00 ;
 reg [31:0] Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 reg [31:0] OOiiILlloiOoI0OlilIOoiiLOOLol0IoI ;
 reg [15:0] OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo ;
 wire [15:0] Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l = (OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo - OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo) ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi <= 16'd0 ;
 O0IILIl0LlliiloOOlliilOilioILILOO <= 16'd0 ;
 OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI <= 16'd0 ;
 OlOO0oILoLOLLLLLllOILOLIilOOLL0oL <= 16'd0 ;
 O0oIIIlIIiOILloLo0lLlILLOL0LIO00O <= 16'd0 ;
 OLLLiliLlOlI00OOlLoLOL00OLoooLIli <= 16'd0 ;
 Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo <= 16'd0 ;
 OIlilLLloioioO00IlooIl0IoOoiOOl0o <= 16'd0 ;
 OLI0O0LOoiLIooi00li0OllLIilLiOiO0 <= 16'd0 ;
 OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO <= 16'd0 ;
 OilloOilLL0Loolo00OIlloliiIoIlOLL <= 16'd0 ;
 O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 <= 16'd0 ;
 O0LoILolI0o00OOoiilOlI0io0O0iiiOi <= 16'd0 ;
 OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol <= 16'd0 ;
 OLlLi0Olo0oloLLoolIi0IIIOlII0LOll <= 16'd0 ;
 OL0OIIiI0loIllilLiIlI0oioI0OloIoL <= 16'd0 ;
 OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil <= 16'd0 ;
 OOI0I0oiooIoOILIL0oLLL0i0iooOL000 <= 16'd0 ;
 O0LL0OoiOLiiII0LooolOliI00oIlIlio <= 16'd0 ;
 O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl <= 16'd0 ;
 OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO <= 16'd0 ;
 OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi <= 16'd0 ;
 OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo <= 16'd0 ;
 OiLOoilOloiOoo0OloLL0llLOIOoLII0O <= 16'd0 ;
 OO0loILiiLolIliIOl0oiloLoioiOLloO <= 16'd0 ;
 OIL0iiOloLOLO0IooOilOiooOilOoLilO <= 16'd0 ;
 OlolILO0OLo0Oi0LiILii00LOlloiLOi0 <= 16'd0 ;
 OL0IoII0L0LLo0IOlLILloi0oi0ilIllI <= 16'd0 ;
 O00OiLOI0i0oL0lOOI0liiol0iLIlOlii <= 16'd0 ;
 O0IoOI0000OlIo0OoiLll0lilIoOLL0ll <= 16'd0 ;
 O0LlIILiOiOioLLoi00lIOi0OI00lOO0I <= 16'd0 ;
 O0LOIioI0oLioOILLLOi0I0IO0ILoioLO <= 16'd0 ;
 end
 else if ( O0oill0llILOilo0i0LIoOLIoolL0Il0o && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] ) OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] && ( OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0]) ) O0IILIl0LlliiloOOlliilOilioILILOO <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1:0]) ) OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2:0]) ) OlOO0oILoLOLLLLLllOILOLIilOOLL0oL <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3:0]) ) O0oIIIlIIiOILloLo0lLlILLOL0LIO00O <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4:0]) ) OLLLiliLlOlI00OOlLoLOL00OLoooLIli <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5:0]) ) Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6:0]) ) OIlilLLloioioO00IlooIl0IoOoiOOl0o <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7:0]) ) OLI0O0LOoiLIooi00li0OllLIilLiOiO0 <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8:0]) ) OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9:0]) ) OilloOilLL0Loolo00OIlloliiIoIlOLL <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10:0]) ) O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11:0]) ) O0LoILolI0o00OOoiilOlI0io0O0iiiOi <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12:0]) ) OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13:0]) ) OLlLi0Olo0oloLLoolIi0IIIOlII0LOll <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14:0]) ) OL0OIIiI0loIllilLiIlI0oioI0OloIoL <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15:0]) ) OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16:0]) ) OOI0I0oiooIoOILIL0oLLL0i0iooOL000 <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17:0]) ) O0LL0OoiOLiiII0LooolOliI00oIlIlio <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18:0]) ) O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19:0]) ) OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20:0]) ) OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21:0]) ) OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22:0]) ) OiLOoilOloiOoo0OloLL0llLOIOoLII0O <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23:0]) ) OO0loILiiLolIliIOl0oiloLoioiOLloO <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24:0]) ) OIL0iiOloLOLO0IooOilOiooOilOoLilO <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25:0]) ) OlolILO0OLo0Oi0LiILii00LOlloiLOi0 <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26:0]) ) OL0IoII0L0LLo0IOlLILloi0oi0ilIllI <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27:0]) ) O00OiLOI0i0oL0lOOI0liiol0iLIlOlii <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28:0]) ) O0IoOI0000OlIo0OoiLll0lilIoOLL0ll <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29:0]) ) O0LlIILiOiOioLLoi00lIOi0OI00lOO0I <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30:0]) ) O0LOIioI0oLioOILLLOi0I0IO0ILoioLO <= OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli ) begin
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ) OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ) O0IILIl0LlliiloOOlliilOilioILILOO <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ) OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ) OlOO0oILoLOLLLLLllOILOLIilOOLL0oL <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ) O0oIIIlIIiOILloLo0lLlILLOL0LIO00O <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ) OLLLiliLlOlI00OOlLoLOL00OLoooLIli <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ) Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ) OIlilLLloioioO00IlooIl0IoOoiOOl0o <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ) OLI0O0LOoiLIooi00li0OllLIilLiOiO0 <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ) OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ) OilloOilLL0Loolo00OIlloliiIoIlOLL <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ) O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ) O0LoILolI0o00OOoiilOlI0io0O0iiiOi <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ) OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ) OLlLi0Olo0oloLLoolIi0IIIOlII0LOll <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ) OL0OIIiI0loIllilLiIlI0oioI0OloIoL <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ) OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ) OOI0I0oiooIoOILIL0oLLL0i0iooOL000 <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ) O0LL0OoiOLiiII0LooolOliI00oIlIlio <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ) O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ) OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ) OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ) OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ) OiLOoilOloiOoo0OloLL0llLOIOoLII0O <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ) OO0loILiiLolIliIOl0oiloLoioiOLloO <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ) OIL0iiOloLOLO0IooOilOiooOilOoLilO <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ) OlolILO0OLo0Oi0LiILii00LOlloiLOi0 <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ) OL0IoII0L0LLo0IOlLILloi0oi0ilIllI <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ) O00OiLOI0i0oL0lOOI0liiol0iLIlOlii <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ) O0IoOI0000OlIo0OoiLll0lilIoOLL0ll <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ) O0LlIILiOiOioLLoi00lIOi0OI00lOO0I <= 16'd8 ;
 if (~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ) O0LOIioI0oLioOILLLOi0I0IO0ILoioLO <= 16'd8 ;
 end
 else if ( (OOLoL0looIOoioIoOooIoLIiIiLiLoiOl ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) ) begin
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0] ) OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi <= OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1] ) O0IILIl0LlliiloOOlliilOilioILILOO <= O0IILIl0LlliiloOOlliilOilioILILOO + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2] ) OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI <= OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3] ) OlOO0oILoLOLLLLLllOILOLIilOOLL0oL <= OlOO0oILoLOLLLLLllOILOLIilOOLL0oL + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4] ) O0oIIIlIIiOILloLo0lLlILLOL0LIO00O <= O0oIIIlIIiOILloLo0lLlILLOL0LIO00O + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5] ) OLLLiliLlOlI00OOlLoLOL00OLoooLIli <= OLLLiliLlOlI00OOlLoLOL00OLoooLIli + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6] ) Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo <= Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7] ) OIlilLLloioioO00IlooIl0IoOoiOOl0o <= OIlilLLloioioO00IlooIl0IoOoiOOl0o + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8] ) OLI0O0LOoiLIooi00li0OllLIilLiOiO0 <= OLI0O0LOoiLIooi00li0OllLIilLiOiO0 + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9] ) OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO <= OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10] ) OilloOilLL0Loolo00OIlloliiIoIlOLL <= OilloOilLL0Loolo00OIlloliiIoIlOLL + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11] ) O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 <= O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12] ) O0LoILolI0o00OOoiilOlI0io0O0iiiOi <= O0LoILolI0o00OOoiilOlI0io0O0iiiOi + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13] ) OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol <= OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14] ) OLlLi0Olo0oloLLoolIi0IIIOlII0LOll <= OLlLi0Olo0oloLLoolIi0IIIOlII0LOll + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15] ) OL0OIIiI0loIllilLiIlI0oioI0OloIoL <= OL0OIIiI0loIllilLiIlI0oioI0OloIoL + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16] ) OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil <= OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17] ) OOI0I0oiooIoOILIL0oLLL0i0iooOL000 <= OOI0I0oiooIoOILIL0oLLL0i0iooOL000 + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18] ) O0LL0OoiOLiiII0LooolOliI00oIlIlio <= O0LL0OoiOLiiII0LooolOliI00oIlIlio + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19] ) O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl <= O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20] ) OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO <= OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21] ) OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi <= OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22] ) OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo <= OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23] ) OiLOoilOloiOoo0OloLL0llLOIOoLII0O <= OiLOoilOloiOoo0OloLL0llLOIOoLII0O + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24] ) OO0loILiiLolIliIOl0oiloLoioiOLloO <= OO0loILiiLolIliIOl0oiloLoioiOLloO + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25] ) OIL0iiOloLOLO0IooOilOiooOilOoLilO <= OIL0iiOloLOLO0IooOilOiooOilOoLilO + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26] ) OlolILO0OLo0Oi0LiILii00LOlloiLOi0 <= OlolILO0OLo0Oi0LiILii00LOlloiLOi0 + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27] ) OL0IoII0L0LLo0IOlLILloi0oi0ilIllI <= OL0IoII0L0LLo0IOlLILloi0oi0ilIllI + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28] ) O00OiLOI0i0oL0lOOI0liiol0iLIlOlii <= O00OiLOI0i0oL0lOOI0liiol0iLIlOlii + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29] ) O0IoOI0000OlIo0OoiLll0lilIoOLL0ll <= O0IoOI0000OlIo0OoiLll0lilIoOLL0ll + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30] ) O0LlIILiOiOioLLoi00lIOi0OI00lOO0I <= O0LlIILiOiOioLLoi00lIOi0OI00lOO0I + 16'd8 ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31] ) O0LOIioI0oLioOILLLOi0I0IO0ILoioLO <= O0LOIioI0oLioOILLLOi0I0IO0ILoioLO + 16'd8 ;
 end
 else if ((OIoIooIolOilIOlooOlOIIOoilLioOIIO ) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl) ) begin
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0] ) OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi <= OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1] ) O0IILIl0LlliiloOOlliilOilioILILOO <= O0IILIl0LlliiloOOlliilOilioILILOO + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2] ) OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI <= OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3] ) OlOO0oILoLOLLLLLllOILOLIilOOLL0oL <= OlOO0oILoLOLLLLLllOILOLIilOOLL0oL + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4] ) O0oIIIlIIiOILloLo0lLlILLOL0LIO00O <= O0oIIIlIIiOILloLo0lLlILLOL0LIO00O + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5] ) OLLLiliLlOlI00OOlLoLOL00OLoooLIli <= OLLLiliLlOlI00OOlLoLOL00OLoooLIli + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6] ) Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo <= Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7] ) OIlilLLloioioO00IlooIl0IoOoiOOl0o <= OIlilLLloioioO00IlooIl0IoOoiOOl0o + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8] ) OLI0O0LOoiLIooi00li0OllLIilLiOiO0 <= OLI0O0LOoiLIooi00li0OllLIilLiOiO0 + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9] ) OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO <= OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10] ) OilloOilLL0Loolo00OIlloliiIoIlOLL <= OilloOilLL0Loolo00OIlloliiIoIlOLL + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11] ) O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 <= O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12] ) O0LoILolI0o00OOoiilOlI0io0O0iiiOi <= O0LoILolI0o00OOoiilOlI0io0O0iiiOi + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13] ) OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol <= OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14] ) OLlLi0Olo0oloLLoolIi0IIIOlII0LOll <= OLlLi0Olo0oloLLoolIi0IIIOlII0LOll + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15] ) OL0OIIiI0loIllilLiIlI0oioI0OloIoL <= OL0OIIiI0loIllilLiIlI0oioI0OloIoL + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16] ) OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil <= OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17] ) OOI0I0oiooIoOILIL0oLLL0i0iooOL000 <= OOI0I0oiooIoOILIL0oLLL0i0iooOL000 + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18] ) O0LL0OoiOLiiII0LooolOliI00oIlIlio <= O0LL0OoiOLiiII0LooolOliI00oIlIlio + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19] ) O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl <= O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20] ) OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO <= OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21] ) OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi <= OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22] ) OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo <= OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23] ) OiLOoilOloiOoo0OloLL0llLOIOoLII0O <= OiLOoilOloiOoo0OloLL0llLOIOoLII0O + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24] ) OO0loILiiLolIliIOl0oiloLoioiOLloO <= OO0loILiiLolIliIOl0oiloLoioiOLloO + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25] ) OIL0iiOloLOLO0IooOilOiooOilOoLilO <= OIL0iiOloLOLO0IooOilOiooOilOoLilO + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26] ) OlolILO0OLo0Oi0LiILii00LOlloiLOi0 <= OlolILO0OLo0Oi0LiILii00LOlloiLOi0 + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27] ) OL0IoII0L0LLo0IOlLILloi0oi0ilIllI <= OL0IoII0L0LLo0IOlLILloi0oi0ilIllI + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28] ) O00OiLOI0i0oL0lOOI0liiol0iLIlOlii <= O00OiLOI0i0oL0lOOI0liiol0iLIlOlii + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29] ) O0IoOI0000OlIo0OoiLll0lilIoOLL0ll <= O0IoOI0000OlIo0OoiLll0lilIoOLL0ll + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30] ) O0LlIILiOiOioLLoi00lIOi0OI00lOO0I <= O0LlIILiOiOioLLoi00lIOi0OI00lOO0I + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 if (OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31] ) O0LOIioI0oLioOILLLOi0I0IO0ILoioLO <= O0LOIioI0oLioOILLLOi0I0IO0ILoioLO + OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= 16'd0 ;
 end
 else if ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI&&OOOLiLOilooIi0Iio00ilILoLIILOoOoI&&(|OI00OiLolooiIIiiILoIliO0O0loolIlI) ) begin
 case (OI00OiLolooiIIiiILoIliO0O0loolIlI) 32'h0000_0001: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OiILoIoLOoilLiOllLIooIL0L0Ooo0iLi ;
 32'h0000_0002: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0IILIl0LlliiloOOlliilOilioILILOO ;
 32'h0000_0004: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OLllIo0il0iOoLIli0iIoIO0iI0Oi0IlI ;
 32'h0000_0008: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OlOO0oILoLOLLLLLllOILOLIilOOLL0oL ;
 32'h0000_0010: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0oIIIlIIiOILloLo0lLlILLOL0LIO00O ;
 32'h0000_0020: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OLLLiliLlOlI00OOlLoLOL00OLoooLIli ;
 32'h0000_0040: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= Oooi0Ol0oLI0L0OOOO0oOILIoOOoiI0Oo ;
 32'h0000_0080: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OIlilLLloioioO00IlooIl0IoOoiOOl0o ;
 32'h0000_0100: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OLI0O0LOoiLIooi00li0OllLIilLiOiO0 ;
 32'h0000_0200: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOLIi0lLOOLILLoOIIOlLOIoioOLloIOO ;
 32'h0000_0400: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OilloOilLL0Loolo00OIlloliiIoIlOLL ;
 32'h0000_0800: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0l0LlO0oLIi0lLoo0IoLli0LoIOLiil0 ;
 32'h0000_1000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0LoILolI0o00OOoiilOlI0io0O0iiiOi ;
 32'h0000_2000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OO0iLoI0oIIi0IOoloOiIo0iIlO0oI0Ol ;
 32'h0000_4000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OLlLi0Olo0oloLLoolIi0IIIOlII0LOll ;
 32'h0000_8000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OL0OIIiI0loIllilLiIlI0oioI0OloIoL ;
 32'h0001_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OoLiIL0I0il0IoOiOlOLO00oIioOo0Iil ;
 32'h0002_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOI0I0oiooIoOILIL0oLLL0i0iooOL000 ;
 32'h0004_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0LL0OoiOLiiII0LooolOliI00oIlIlio ;
 32'h0008_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0IoLiOIOIlIo0iIlOLIioiLI0LOIIiOl ;
 32'h0010_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOl0LLiOiIoiOIlllL0oiLiLooLOioiLO ;
 32'h0020_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OIIO00iLLlILOLOooIOOOLLi0IiOOIOIi ;
 32'h0040_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OLlOL0oI0OLOI0IlLloLoiIIioLLOL0Oo ;
 32'h0080_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OiLOoilOloiOoo0OloLL0llLOIOoLII0O ;
 32'h0100_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OO0loILiiLolIliIOl0oiloLoioiOLloO ;
 32'h0200_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OIL0iiOloLOLO0IooOilOiooOilOoLilO ;
 32'h0400_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OlolILO0OLo0Oi0LiILii00LOlloiLOi0 ;
 32'h0800_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OL0IoII0L0LLo0IOlLILloi0oi0ilIllI ;
 32'h1000_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O00OiLOI0i0oL0lOOI0liiol0iLIlOlii ;
 32'h2000_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0IoOI0000OlIo0OoiLll0lilIoOLL0ll ;
 32'h4000_0000: OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0LlIILiOiOioLLoi00lIOi0OI00lOO0I ;
 default : OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= O0LOIioI0oLioOILLLOi0I0IO0ILoioLO ;
 endcase end
 else if (OiL0LolLLIOlliloII00llOil0oIlOiIo && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=16'd8) ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo + 16'd8 ;
 end
 else if (O0llIOIliLOO0iiOoO0OO0lIOloLoII0I && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l) ) begin
 OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo <= OOoi0IIoiILOiOLIOo0LiOl0lOoLOL0Lo + Oii0ILIlIiIIiiIOI0OLillOolIIoOO0l ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= 16'd0 ;
 end
 else if ( |OI00OiLolooiIIiiILoIliO0O0loolIlI ) begin
 case (OI00OiLolooiIIiiILoIliO0O0loolIlI) 32'h0000_0001: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OlOiLoIOLoOOiOLiOoOL0iOloioliL0OI ;
 32'h0000_0002: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OOL0LOOi0lL0Ooo0ooOLLLOO0OLo0iolL ;
 32'h0000_0004: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= Oo0OiL0Lll000LlioLiooLOLloiLiliii ;
 32'h0000_0008: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OIoOlOlloI0oio0LLOIOIlOoOOlIoOLoI ;
 32'h0000_0010: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OioiIooIlil0liIiOIi0lLLIllOioioli ;
 32'h0000_0020: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OL0OlLIiiOl00iL0LIOo0LiIlOIOO0II0 ;
 32'h0000_0040: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OlLloLOlOi0iIiLIlOlLio000LLOLILli ;
 32'h0000_0080: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OIio0oi0oL0l0llO0ii0lILOio0OOl0I0 ;
 32'h0000_0100: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OOlILOLoilIOloioiIoOLI0L0ooLO0Lll ;
 32'h0000_0200: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OolOlIOiIIoII0ll0IllLoOiIllIilOoO ;
 32'h0000_0400: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OOIiiol0IOILiLloOLiLOIIlIIolooOIO ;
 32'h0000_0800: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OiLi0I0LLio0iioLOi0OlLl0l0OLioIoO ;
 32'h0000_1000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OILili00ILILlO0LIoLlll0oliLio0liL ;
 32'h0000_2000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OoILoooiioLLiIIIoiIoiOIO0OllIlIlL ;
 32'h0000_4000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OiOILIIOL0OI0lIIoIooiO0ioLOIII0lO ;
 32'h0000_8000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OIiiiIlLolLIoIioOoOolloi0L0loLoIL ;
 32'h0001_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OILO0OL0LOIiIIoiiOLIIo00ol0IIoloO ;
 32'h0002_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= O0oLLIlOIlOiiLiloo0OoO0Liio0OL0II ;
 32'h0004_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OIOIO0L00OiLLOLLiOo0IliI0OOOoIIoO ;
 32'h0008_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OOlO0o0i0Io0IOllLoIloiioiliOOlIII ;
 32'h0010_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OLI00ioL0IlLOOlIoillOoOIoLiOLIi0I ;
 32'h0020_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= O0OliLI0l00IIl0oi0ioOOiiLLOL0oLi0 ;
 32'h0040_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OlOlLO00i0Oiooo0lLollo0IILIlLO0OI ;
 32'h0080_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OLLliI0IiOiollllIOOLL0oL0IlllO0oI ;
 32'h0100_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OLO00iLliol0LLIOOIIO0IiLIllO0IL0O ;
 32'h0200_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= O0OII0Ili0ilol00OLOLoiOl0OlLo0liO ;
 32'h0400_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OOL0lolilI0oIloIoIIILooo0lOLOlolI ;
 32'h0800_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OlIo0o0iI0lOOiiOIoO0OOOoliOLoL0ll ;
 32'h1000_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OIO00IOolLoOoOL0ILI00i0olI0IiiOOo ;
 32'h2000_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OI0LoiOlOOO0ooL00IiLLoi00IOIl0llO ;
 32'h4000_0000: OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OLlOOlIoLlo0iiooIIlllO0ooloL0iIi0 ;
 default : OiO0iOlio0Ii0liiOIO0OLIiL000oIIoo <= OIoiIlOo00oL0iL0o0iooollLlilLoIIo ;
 endcase end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0OlOIIOOIOIioo00liool0iIiI0I0Lll <= 1'd0 ;
 O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii <= 4'd0 ;
 OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l <= 1'd0 ;
 OIiOIl0O0OLllloOl0oOoLoIllIL0illO <= 1'd0 ;
 Oi0loi0OllIlIoI0ILloIllILIO0IIo0I <= 64'd0 ;
 OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i <= 16'd0 ;
 OOloOOOOiILOioIlIOO0oILilOLLL00OO <= 16'd0 ;
 OOIlIOO0IL0OoLli0IoliIioOOlIILlii <= 32'd0 ;
 OioOlll0OooLLL0IIIIIli0ollooo0L0L <= 1'd0 ;
 OooOLOOliIlIOlio00OO0oloLoOi0lliO <= 32'd0 ;
 OoI0IoiILOOLILioiioIOoOLioiiOlIio <= 1'd0 ;
 OoLOIol0OLIIiloO0oLoiliOl0LilIolI <= 'd0 ;
 end
 else begin
 O0OlOIIOOIOIioo00liool0iIiI0I0Lll <= OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii <= OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII : O0Ll0OO0LLOIiiLiiOlloolOOIolLLIii ;
 OOLOoIoI0lO0OI0iioOOo0oiOlIOILO0l <= OOLOoolOi0LIo0olO0loLllIlllIiiIiI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 OIiOIl0O0OLllloOl0oOoLoIllIL0illO <= OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 Oi0loi0OllIlIoI0ILloIllILIO0IIo0I <= OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? OLLOooI0ILL00ILloiliILLLiioooLliI : Oi0loi0OllIlIoI0ILloIllILIO0IIo0I ;
 OoLOIol0OLIIiloO0oLoiliOl0LilIolI <= OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? OILoli0OIOIIOI0OiliOo0i0OLoliOOiI : OoLOIol0OLIIiloO0oLoiliOl0LilIolI ;
 OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i <= OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI : OIllLOoiL0IIoiOooLOlLoLoi0O0lIO0i ;
 OOloOOOOiILOioIlIOO0oILilOLLL00OO <= OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? OilOOioILlOIIOL0iioIOIi0oloooOoLl : OOloOOOOiILOioIlIOO0oILilOLLL00OO ;
 OOIlIOO0IL0OoLli0IoliIioOOlIILlii <= OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? OI00OiLolooiIIiiILoIliO0O0loolIlI : OOIlIOO0IL0OoLli0IoliIioOOlIILlii ;
 OioOlll0OooLLL0IIIIIli0ollooo0L0L <= OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? (|OI00OiLolooiIIiiILoIliO0O0loolIlI) : OioOlll0OooLLL0IIIIIli0ollooo0L0L ;
 OooOLOOliIlIOlio00OO0oloLoOi0lliO <= OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? OIIOLLOIlOlLoi0oiOioLilOiioiiliLO : OooOLOOliIlIOlio00OO0oloLoOi0lliO ;
 OoI0IoiILOOLILioiioIOoOLioiiOlIio <= OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && OOOLiLOilooIi0Iio00ilILoLIILOoOoI ? (|OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo) : OoI0IoiILOOLILioiioIOoOLioiiOlIio ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI <= 32'd0 ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli && (OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ;
 end
 else if (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli && (|OolIOLOooiLLIllI0LOLIolllLoilolIl) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8 ) ) begin
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 0] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 1] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 2] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 3] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 4] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 5] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 6] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 7] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 8] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[ 9] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[10] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[11] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[12] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[13] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[14] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[15] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[16] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[17] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[18] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[19] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[20] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[21] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[22] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[23] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[24] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[25] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[26] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[27] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[28] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[29] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[30] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ;
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI[31] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ;
 end
 else if (Oi0OIIIIi0I0iIlOIIIlollIi0iOoOIII) begin
 OOiiILlloiOoI0OlilIOoiiLOOLol0IoI <= 32'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O <= 32'd0 ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli && (OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 0] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 1] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 2] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 3] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 4] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 5] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 6] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 7] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 8] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 9] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[10] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[11] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[12] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[13] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[14] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[15] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[16] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[17] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[18] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[19] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[20] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[21] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[22] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[23] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[24] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[25] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[26] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[27] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[28] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[29] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[30] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[31] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ;
 end
 else if (OI0o0L00o0ilL0ioLLlLO0i0oIilolOIL && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli && (|OolIOLOooiLLIllI0LOLIolllLoilolIl) && (OolIOLOooiLLIllI0LOLIolllLoilolIl<=16'd8 ) ) begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 0] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 1] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 2] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 3] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 4] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 5] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 6] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 7] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 8] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 9] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[10] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[11] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[12] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[13] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[14] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[15] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[16] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[17] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[18] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[19] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[20] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[21] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[22] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[23] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[24] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[25] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[26] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[27] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[28] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[29] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[30] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29:0]) ;
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[31] <= ~OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && (&OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30:0]) ;
 end
 else begin
 OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O <= 32'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OLOoliOOlOIIIioiilio0liLil0o0I000 <= 32'd0 ;
 end
 else if ( OlliILlLOilOl0LO0O0OilooiIIiOi0Ll && (OolIOLOooiLLIllI0LOLIolllLoilolIl<(O0OiLI0oloiOLoi0lOlo0oLOOilLooLLo+16'd4)) && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=6'd8) && OI0OOoIliioLOLiI0IOOiL0l0o0OiOIo0 && O0Loo0iiI0OlLOlOIiILOooOOlIoioOli && (OILIloOoilLIL00IIOoOilLOO0L0iiIOO==16'h0200)&&(O0oLLi0Ill00l0lioiLioiooIllloIiIl==32'h0100_044c) ) begin
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 0] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 1] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] && ( OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 2] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 3] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 4] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 5] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 6] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 7] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 8] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 9] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[10] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[11] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[12] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[13] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[14] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[15] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[16] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[17] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[18] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[19] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[20] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[21] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[22] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[23] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[24] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[25] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[26] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[27] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[28] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[29] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[30] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[31] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30:0]) ;
 end
 else if ( O0oill0llILOilo0i0LIoOLIoolL0Il0o && (O0IOooLliOlIllOliILoolIIoIiO0Ilol>=OolIOLOooiLLIllI0LOLIolllLoilolIl ) ) begin
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 0] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 1] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] && ( OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 2] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 3] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 4] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 5] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 6] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 7] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 8] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[ 9] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[10] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[11] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[12] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[13] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[14] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[15] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[16] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[17] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[18] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[19] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[20] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[21] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[22] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[23] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[24] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[25] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[26] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[27] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[28] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[29] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[30] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29:0]) ;
 OLOoliOOlOIIIioiilio0liLil0o0I000[31] <= ~OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] && (&OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30:0]) ;
 end
 else begin
 OLOoliOOlOIIIioiilio0liLil0o0I000 <= 32'd0 ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI <= 32'd0 ;
 end
 else if ( |OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ) begin
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 0] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 1] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 2] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 3] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 4] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 5] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 6] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 7] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 8] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 9] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[10] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[11] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[12] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[13] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[14] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[15] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[16] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[17] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[18] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[19] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[20] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[21] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[22] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[23] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[24] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[25] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[26] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[27] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[28] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[29] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[30] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] <= OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[31] ? 1'd1 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] ;
 end
 else if ( |OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ) begin
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 0] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 1] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 2] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 3] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 4] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 5] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 6] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 7] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 8] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 9] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[10] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[11] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[12] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[13] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[14] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[15] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[16] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[17] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[18] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[19] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[20] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[21] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[22] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[23] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[24] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[25] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[26] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[27] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[28] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[29] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[30] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[31] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] ;
 end
 else if ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && (|OI00OiLolooiIIiiILoIliO0O0loolIlI) ) begin
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 0] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 1] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 2] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 3] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 4] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 5] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 6] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 7] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 8] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 9] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[10] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[11] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[12] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[13] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[14] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[15] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[16] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[17] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[18] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[19] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[20] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[21] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[22] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[23] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[24] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[25] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[26] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[27] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[28] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[29] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[30] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] ;
 OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[31] ? 1'd0 : OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO <= 32'd0 ;
 end
 else if ( |OLOoliOOlOIIIioiilio0liLil0o0I000 ) begin
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 0] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 1] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 2] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 3] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 4] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 5] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 6] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 7] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 8] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] <= OLOoliOOlOIIIioiilio0liLil0o0I000[ 9] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] <= OLOoliOOlOIIIioiilio0liLil0o0I000[10] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] <= OLOoliOOlOIIIioiilio0liLil0o0I000[11] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] <= OLOoliOOlOIIIioiilio0liLil0o0I000[12] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] <= OLOoliOOlOIIIioiilio0liLil0o0I000[13] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] <= OLOoliOOlOIIIioiilio0liLil0o0I000[14] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] <= OLOoliOOlOIIIioiilio0liLil0o0I000[15] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] <= OLOoliOOlOIIIioiilio0liLil0o0I000[16] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] <= OLOoliOOlOIIIioiilio0liLil0o0I000[17] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] <= OLOoliOOlOIIIioiilio0liLil0o0I000[18] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] <= OLOoliOOlOIIIioiilio0liLil0o0I000[19] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] <= OLOoliOOlOIIIioiilio0liLil0o0I000[20] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] <= OLOoliOOlOIIIioiilio0liLil0o0I000[21] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] <= OLOoliOOlOIIIioiilio0liLil0o0I000[22] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] <= OLOoliOOlOIIIioiilio0liLil0o0I000[23] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] <= OLOoliOOlOIIIioiilio0liLil0o0I000[24] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] <= OLOoliOOlOIIIioiilio0liLil0o0I000[25] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] <= OLOoliOOlOIIIioiilio0liLil0o0I000[26] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] <= OLOoliOOlOIIIioiilio0liLil0o0I000[27] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] <= OLOoliOOlOIIIioiilio0liLil0o0I000[28] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] <= OLOoliOOlOIIIioiilio0liLil0o0I000[29] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] <= OLOoliOOlOIIIioiilio0liLil0o0I000[30] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] <= OLOoliOOlOIIIioiilio0liLil0o0I000[31] ? 1'd1 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] ;
 end
 else if ( |OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ) begin
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 0] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 1] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 2] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 3] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 4] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 5] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 6] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 7] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 8] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[ 9] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[10] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[11] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[12] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[13] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[14] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[15] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[16] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[17] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[18] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[19] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[20] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[21] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[22] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[23] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[24] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[25] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[26] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[27] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[28] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[29] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[30] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] <= OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI[31] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] ;
 end
 else if ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI && (|OI00OiLolooiIIiiILoIliO0O0loolIlI) ) begin
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 0] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 0] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 1] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 1] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 2] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 2] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 3] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 3] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 4] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 4] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 5] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 5] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 6] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 6] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 7] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 7] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 8] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 8] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[ 9] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[ 9] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[10] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[10] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[11] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[11] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[12] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[12] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[13] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[13] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[14] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[14] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[15] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[15] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[16] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[16] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[17] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[17] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[18] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[18] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[19] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[19] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[20] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[20] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[21] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[21] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[22] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[22] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[23] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[23] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[24] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[24] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[25] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[25] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[26] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[26] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[27] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[27] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[28] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[28] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[29] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[29] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[30] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[30] ;
 OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] <= OI00OiLolooiIIiiILoIliO0O0loolIlI[31] ? 1'd0 : OioL00ILO0li0IO0LIlIO00lL0I0OllIO[31] ;
 end
 end
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OliiILooLoLLIi0IliLO0OO0OOiololoL <= 32'd0 ;
 Oll0lolIi00IiOOiIl00OI0OLoIioOLOl <= 32'd0 ;
 OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I <= 32'd0 ;
 OOOiOlOLli0LLiOOLILIllil0OiLLli0L <= 32'd0 ;
 O0LiLoL0IooiOILoioILLLLli00o0LI0I <= 32'd0 ;
 OIolIiLOiOLoO00oiliiollllO0l0OloO <= 32'd0 ;
 Oil0OiILooLiiioloiiI0oLLlOlLllo0i <= 32'd0 ;
 OI0LoL000LIII0lI0LL0LoilIiIlLLiOl <= 32'd0 ;
 OoiLi0oolILIllloliLiL0LolIliiLOlo <= 32'd0 ;
 OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO <= 32'd0 ;
 OioooOOI00ollOl0LiLIl0LIliO00OOii <= 32'd0 ;
 OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl <= 32'd0 ;
 OoolIOILLooLiOLlLiIoO00OooLLL0LLO <= 32'd0 ;
 OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0 <= 32'd0 ;
 OoIIliiLlI0OilooiiILLLOL0oII0ILio <= 32'd0 ;
 OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i <= 32'd0 ;
 OliilLooOIL0lio0OOioLLoLoLOlioIio <= 32'd0 ;
 OolioiLoIlIlolO0ooiO0OLOoIlIllIi0 <= 32'd0 ;
 OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo <= 32'd0 ;
 OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo <= 32'd0 ;
 O0iiOolLIl0iOLOiLOOLII00IloOo0li0 <= 32'd0 ;
 OLilOOlILoL0oioOOOlOLlOl0li0lIli0 <= 32'd0 ;
 OlIIiOliliiioo0LO0I0IIOIiLLooI0lI <= 32'd0 ;
 OiOllilOOiI0II0IIilo0IllOOIIIoLii <= 32'd0 ;
 OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI <= 32'd0 ;
 OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l <= 32'd0 ;
 OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0 <= 32'd0 ;
 OloOLL0I00I0oIIILLo0Ol0Il0lIILL00 <= 32'd0 ;
 OioiIOLioLOlOoliOlLli0i0IolIlOLiL <= 32'd0 ;
 OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI <= 32'd0 ;
 OiIooILlOili0io0LiiiILIloOi0lIIOl <= 32'd0 ;
 OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00 <= 32'd0 ;
 end
 else if ( |OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ) begin
 OliiILooLoLLIi0IliLO0OO0OOiololoL <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 0]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OliiILooLoLLIi0IliLO0OO0OOiololoL ;
 Oll0lolIi00IiOOiIl00OI0OLoIioOLOl <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 1]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : Oll0lolIi00IiOOiIl00OI0OLoIioOLOl ;
 OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 2]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I ;
 OOOiOlOLli0LLiOOLILIllil0OiLLli0L <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 3]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OOOiOlOLli0LLiOOLILIllil0OiLLli0L ;
 O0LiLoL0IooiOILoioILLLLli00o0LI0I <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 4]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : O0LiLoL0IooiOILoioILLLLli00o0LI0I ;
 OIolIiLOiOLoO00oiliiollllO0l0OloO <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 5]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OIolIiLOiOLoO00oiliiollllO0l0OloO ;
 Oil0OiILooLiiioloiiI0oLLlOlLllo0i <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 6]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : Oil0OiILooLiiioloiiI0oLLlOlLllo0i ;
 OI0LoL000LIII0lI0LL0LoilIiIlLLiOl <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 7]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OI0LoL000LIII0lI0LL0LoilIiIlLLiOl ;
 OoiLi0oolILIllloliLiL0LolIliiLOlo <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 8]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OoiLi0oolILIllloliLiL0LolIliiLOlo ;
 OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[ 9]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO ;
 OioooOOI00ollOl0LiLIl0LIliO00OOii <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[10]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OioooOOI00ollOl0LiLIl0LIliO00OOii ;
 OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[11]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl ;
 OoolIOILLooLiOLlLiIoO00OooLLL0LLO <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[12]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OoolIOILLooLiOLlLiIoO00OooLLL0LLO ;
 OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[13]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0 ;
 OoIIliiLlI0OilooiiILLLOL0oII0ILio <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[14]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OoIIliiLlI0OilooiiILLLOL0oII0ILio ;
 OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[15]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i ;
 OliilLooOIL0lio0OOioLLoLoLOlioIio <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[16]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OliilLooOIL0lio0OOioLLoLoLOlioIio ;
 OolioiLoIlIlolO0ooiO0OLOoIlIllIi0 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[17]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OolioiLoIlIlolO0ooiO0OLOoIlIllIi0 ;
 OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[18]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo ;
 OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[19]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo ;
 O0iiOolLIl0iOLOiLOOLII00IloOo0li0 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[20]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : O0iiOolLIl0iOLOiLOOLII00IloOo0li0 ;
 OLilOOlILoL0oioOOOlOLlOl0li0lIli0 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[21]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OLilOOlILoL0oioOOOlOLlOl0li0lIli0 ;
 OlIIiOliliiioo0LO0I0IIOIiLLooI0lI <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[22]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OlIIiOliliiioo0LO0I0IIOIiLLooI0lI ;
 OiOllilOOiI0II0IIilo0IllOOIIIoLii <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[23]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OiOllilOOiI0II0IIilo0IllOOIIIoLii ;
 OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[24]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI ;
 OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[25]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l ;
 OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[26]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0 ;
 OloOLL0I00I0oIIILLo0Ol0Il0lIILL00 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[27]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OloOLL0I00I0oIIILLo0Ol0Il0lIILL00 ;
 OioiIOLioLOlOoliOlLli0i0IolIlOLiL <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[28]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OioiIOLioLOlOoliOlLli0i0IolIlOLiL ;
 OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[29]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI ;
 OiIooILlOili0io0LiiiILIloOi0lIIOl <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[30]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OiIooILlOili0io0LiiiILIloOi0lIIOl ;
 OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00 <= (OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O[31]) ? OO0liOO0iOOIioool0OoLliiiI0l0ilOo + 1'd1 : OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00 ;
 end
 end
 reg OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= 32'd0 ;
 OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl <= 1'd0 ;
 end
 else begin
 OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl <= |Oo0LLillol0loLIo0iOl0oOLlIOlILoIO ;
 case (Oo0LLillol0loLIo0iOl0oOLlIOlILoIO) 32'h0000_0001: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLl0loOLioi0II0ioOi0iLIi0iLIOIOlO) ;
 32'h0000_0002: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLlOiiLlLoolliOiO0i0lOloio0L0oL00) ;
 32'h0000_0004: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OilOI0i0lloo0Lll000I0OIoIOI0lioiO) ;
 32'h0000_0008: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlooiiLooL0L00oIIiioLloiIolOoOlLo) ;
 32'h0000_0010: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLo0LOlILllLILOIiiiL0LIlLIoLlO0II) ;
 32'h0000_0020: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OiiOioOIO00LOOLilooiooo0olO0illo0) ;
 32'h0000_0040: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLl0LoLoii00oiOOoilollii000iIOlOI) ;
 32'h0000_0080: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLlil0000Oiil0IOOLiloIlliOoLLol0L) ;
 32'h0000_0100: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OIOl0liIiI0OLOIO0L0OLilIi0iILI0oI) ;
 32'h0000_0200: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OO0OOILiO000LOILL0OllLi0l0oliLOo0) ;
 32'h0000_0400: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLiLllIIIlo0llILiLloLOoooOLOilI0l) ;
 32'h0000_0800: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (Oo0L0IOLoOill0ilOIi0IOiiooLLIOLIl) ;
 32'h0000_1000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OiL0IiiliiioOOLliLiiLILlIOloOLL0L) ;
 32'h0000_2000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlIi0ili0IIo0Oi00OLOOLLioOL0lLIOi) ;
 32'h0000_4000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OllLOLiIilI0oili000OiLilLioIOoIl0) ;
 32'h0000_8000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOooI0loOL0iiOIoOili0OOOLLiiIiLOl) ;
 32'h0001_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OLIIiIIIOILl0loi0lO0IiOoolLIloi00) ;
 32'h0002_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OoOillIILLoLoOioLloli0OLILlIOOoLo) ;
 32'h0004_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlOlO00LLloOiOolOiOLOIiloLil0L0LI) ;
 32'h0008_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OooL0I0IiIOOiLLOiLIII0oIiLlIOiloO) ;
 32'h0010_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlOLIILoL0ll0oooOo0OIoLoOoiLIolol) ;
 32'h0020_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OIlLOILiLLo0ol0OLlI0IILilILLLlILO) ;
 32'h0040_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (O0OL0LiIIIlIiOOIoOOoI0IIoIoOiI00i) ;
 32'h0080_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (Oo0l0OL0OliIlIIIllo0IliIO0O0LlllL) ;
 32'h0100_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOiIlillllLOI0oOOoILlol0ILoIoOLil) ;
 32'h0200_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOIiO0olO0OLlo0liIoiOioiIO00oOIiL) ;
 32'h0400_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (O0Illi0IOIoiO0I0IiLLIo0ilLiOOILi0) ;
 32'h0800_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OOLoILl00II0l0O0LiIOOo0Oiiii0oo0l) ;
 32'h1000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlolLlliLo0O0l0lOOolL0ioI0O0Li00l) ;
 32'h2000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (Oo0oI0oLOLlloloiiLIIol0LilOlOIliI) ;
 32'h4000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OlLOOOOlliLoi0IiLOoLL0iiloiOLOLoo) ;
 32'h8000_0000: Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= (OoiLlL0oiiIloLOoloIL0oLii00IIIoII) ;
 default : Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO <= Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO ;
 endcase end
 end
 reg [1:0] OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO ;
 reg [1:0] OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i ;
 reg [1:0] OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo ;
 reg [1:0] OiLoOlOLii00LILIoloiioLiIoIoioO0L ;
 reg [1:0] O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I ;
 reg [1:0] OIoLLIoLLLIILi0oi00LolIolIIoliiiI ;
 reg [1:0] Oi0OollLl0olLol00i0iOOLI0ILliIIIi ;
 reg [1:0] OO0Ii0IOoilLoILLOIIli0LOLilliLOlI ;
 reg [1:0] O0llOO0ilOIiiioOi0Oloo0IlIILOIlio ;
 reg [1:0] Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo ;
 reg [1:0] O0Iliiill00LoolO00Oo0oI00OoolLlLo ;
 reg [1:0] O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI ;
 reg [1:0] OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O ;
 reg [1:0] OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo ;
 reg [1:0] OoILiLOioiOIolLloILoIOLio0iLLoiii ;
 reg [1:0] OLoO0iLi00loILiIo0OlOolilIilOlIii ;
 reg [1:0] OIIoO0IiLililLIoiilIl00olLoOIlLoL ;
 reg [1:0] OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo ;
 reg [1:0] OIoI0IOlOLiOllo0iooll00o0lOOoIooo ;
 reg [1:0] OOLoioilOIOlOOI0iiII0IIOIL0olIL0O ;
 reg [1:0] OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL ;
 reg [1:0] OIIi0OoOILoL0LLlLiIOILill0o0ll0OI ;
 reg [1:0] OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo ;
 reg [1:0] OLoiILloilO0IIiOOlLoo0LL0ILllliLO ;
 reg [1:0] OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L ;
 reg [1:0] OILlI00OIL0i0OOl0IlOoloII0o0oOlOL ;
 reg [1:0] OlLIlilLII00OliliLLiLIII0000Ll0o0 ;
 reg [1:0] OooIIILiI0ILoOlO0o0il0LiOoLLLILiO ;
 reg [1:0] OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI ;
 reg [1:0] OlL0O0LOLillLLIOoOLl0lOOioOiliOol ;
 reg [1:0] OilIIlLl0oo0iilIiiOlilILOlo0IIOOI ;
 reg [1:0] OOI0IILoliiOO0lioiOiO0iloIiOlIlL0 ;
 always@ ( negedge OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI or posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if (~OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 O0I0oI0I000LllOOI0L0lOlIl000LIioO <= 32'd0 ;
 OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO <= 2'd0 ;
 OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i <= 2'd0 ;
 OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo <= 2'd0 ;
 OiLoOlOLii00LILIoloiioLiIoIoioO0L <= 2'd0 ;
 O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I <= 2'd0 ;
 OIoLLIoLLLIILi0oi00LolIolIIoliiiI <= 2'd0 ;
 Oi0OollLl0olLol00i0iOOLI0ILliIIIi <= 2'd0 ;
 OO0Ii0IOoilLoILLOIIli0LOLilliLOlI <= 2'd0 ;
 O0llOO0ilOIiiioOi0Oloo0IlIILOIlio <= 2'd0 ;
 Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo <= 2'd0 ;
 O0Iliiill00LoolO00Oo0oI00OoolLlLo <= 2'd0 ;
 O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI <= 2'd0 ;
 OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O <= 2'd0 ;
 OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo <= 2'd0 ;
 OoILiLOioiOIolLloILoIOLio0iLLoiii <= 2'd0 ;
 OLoO0iLi00loILiIo0OlOolilIilOlIii <= 2'd0 ;
 OIIoO0IiLililLIoiilIl00olLoOIlLoL <= 2'd0 ;
 OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo <= 2'd0 ;
 OIoI0IOlOLiOllo0iooll00o0lOOoIooo <= 2'd0 ;
 OOLoioilOIOlOOI0iiII0IIOIL0olIL0O <= 2'd0 ;
 OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL <= 2'd0 ;
 OIIi0OoOILoL0LLlLiIOILill0o0ll0OI <= 2'd0 ;
 OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo <= 2'd0 ;
 OLoiILloilO0IIiOOlLoo0LL0ILllliLO <= 2'd0 ;
 OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L <= 2'd0 ;
 OILlI00OIL0i0OOl0IlOoloII0o0oOlOL <= 2'd0 ;
 OlLIlilLII00OliliLLiLIII0000Ll0o0 <= 2'd0 ;
 OooIIILiI0ILoOlO0o0il0LiOoLLLILiO <= 2'd0 ;
 OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI <= 2'd0 ;
 OlL0O0LOLillLLIOoOLl0lOOioOiliOol <= 2'd0 ;
 OilIIlLl0oo0iilIiiOlilILOlo0IIOOI <= 2'd0 ;
 OOI0IILoliiOO0lioiOiO0iloIiOlIlL0 <= 2'd0 ;
 end
 else if (OOLOlOo0000iOi0OLOolloLo0iL0iooIi) begin
 O0I0oI0I000LllOOI0L0lOlIl000LIioO <= 32'h0000_0000 ;
 OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO <= 2'd0 ;
 OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i <= 2'd0 ;
 OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo <= 2'd0 ;
 OiLoOlOLii00LILIoloiioLiIoIoioO0L <= 2'd0 ;
 O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I <= 2'd0 ;
 OIoLLIoLLLIILi0oi00LolIolIIoliiiI <= 2'd0 ;
 Oi0OollLl0olLol00i0iOOLI0ILliIIIi <= 2'd0 ;
 OO0Ii0IOoilLoILLOIIli0LOLilliLOlI <= 2'd0 ;
 O0llOO0ilOIiiioOi0Oloo0IlIILOIlio <= 2'd0 ;
 Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo <= 2'd0 ;
 O0Iliiill00LoolO00Oo0oI00OoolLlLo <= 2'd0 ;
 O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI <= 2'd0 ;
 OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O <= 2'd0 ;
 OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo <= 2'd0 ;
 OoILiLOioiOIolLloILoIOLio0iLLoiii <= 2'd0 ;
 OLoO0iLi00loILiIo0OlOolilIilOlIii <= 2'd0 ;
 OIIoO0IiLililLIoiilIl00olLoOIlLoL <= 2'd0 ;
 OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo <= 2'd0 ;
 OIoI0IOlOLiOllo0iooll00o0lOOoIooo <= 2'd0 ;
 OOLoioilOIOlOOI0iiII0IIOIL0olIL0O <= 2'd0 ;
 OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL <= 2'd0 ;
 OIIi0OoOILoL0LLlLiIOILill0o0ll0OI <= 2'd0 ;
 OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo <= 2'd0 ;
 OLoiILloilO0IIiOOlLoo0LL0ILllliLO <= 2'd0 ;
 OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L <= 2'd0 ;
 OILlI00OIL0i0OOl0IlOoloII0o0oOlOL <= 2'd0 ;
 OlLIlilLII00OliliLLiLIII0000Ll0o0 <= 2'd0 ;
 OooIIILiI0ILoOlO0o0il0LiOoLLLILiO <= 2'd0 ;
 OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI <= 2'd0 ;
 OlL0O0LOLillLLIOoOLl0lOOioOiliOol <= 2'd0 ;
 OilIIlLl0oo0iilIiiOlilILOlo0IIOOI <= 2'd0 ;
 OOI0IILoliiOO0lioiOiO0iloIiOlIlL0 <= 2'd0 ;
 end
 else if ( OLoLlLiOlolOil0OLlliIli0Ol0LIOiIl ) begin
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 0] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] && ( (OliiILooLoLLIi0IliLO0OO0OOiololoL==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OliiILooLoLLIi0IliLO0OO0OOiololoL<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 1] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && ( (Oll0lolIi00IiOOiIl00OI0OLoIioOLOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (Oll0lolIi00IiOOiIl00OI0OLoIioOLOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 2] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && ( (OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 3] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && ( (OOOiOlOLli0LLiOOLILIllil0OiLLli0L==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OOOiOlOLli0LLiOOLILIllil0OiLLli0L<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OiLoOlOLii00LILIoloiioLiIoIoioO0L>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 4] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && ( (O0LiLoL0IooiOILoioILLLLli00o0LI0I==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (O0LiLoL0IooiOILoioILLLLli00o0LI0I<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 5] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && ( (OIolIiLOiOLoO00oiliiollllO0l0OloO==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OIolIiLOiOLoO00oiliiollllO0l0OloO<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OIoLLIoLLLIILi0oi00LolIolIIoliiiI>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 6] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && ( (Oil0OiILooLiiioloiiI0oLLlOlLllo0i==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (Oil0OiILooLiiioloiiI0oLLlOlLllo0i<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (Oi0OollLl0olLol00i0iOOLI0ILliIIIi>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 7] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && ( (OI0LoL000LIII0lI0LL0LoilIiIlLLiOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OI0LoL000LIII0lI0LL0LoilIiIlLLiOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OO0Ii0IOoilLoILLOIIli0LOLilliLOlI>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 8] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && ( (OoiLi0oolILIllloliLiL0LolIliiLOlo==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OoiLi0oolILIllloliLiL0LolIliiLOlo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (O0llOO0ilOIiiioOi0Oloo0IlIILOIlio>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 9] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && ( (OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[10] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && ( (OioooOOI00ollOl0LiLIl0LIliO00OOii==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OioooOOI00ollOl0LiLIl0LIliO00OOii<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (O0Iliiill00LoolO00Oo0oI00OoolLlLo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[11] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && ( (OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[12] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && ( (OoolIOILLooLiOLlLiIoO00OooLLL0LLO==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OoolIOILLooLiOLlLiIoO00OooLLL0LLO<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[13] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && ( (OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[14] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && ( (OoIIliiLlI0OilooiiILLLOL0oII0ILio==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OoIIliiLlI0OilooiiILLLOL0oII0ILio<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OoILiLOioiOIolLloILoIOLio0iLLoiii>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[15] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && ( (OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OLoO0iLi00loILiIo0OlOolilIilOlIii>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[16] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && ( (OliilLooOIL0lio0OOioLLoLoLOlioIio==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OliilLooOIL0lio0OOioLLoLoLOlioIio<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OIIoO0IiLililLIoiilIl00olLoOIlLoL>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[17] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && ( (OolioiLoIlIlolO0ooiO0OLOoIlIllIi0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OolioiLoIlIlolO0ooiO0OLOoIlIllIi0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[18] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && ( (OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OIoI0IOlOLiOllo0iooll00o0lOOoIooo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[19] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && ( (OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OOLoioilOIOlOOI0iiII0IIOIL0olIL0O>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[20] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && ( (O0iiOolLIl0iOLOiLOOLII00IloOo0li0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (O0iiOolLIl0iOLOiLOOLII00IloOo0li0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[21] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && ( (OLilOOlILoL0oioOOOlOLlOl0li0lIli0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OLilOOlILoL0oioOOOlOLlOl0li0lIli0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OIIi0OoOILoL0LLlLiIOILill0o0ll0OI>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[22] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && ( (OlIIiOliliiioo0LO0I0IIOIiLLooI0lI==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OlIIiOliliiioo0LO0I0IIOIiLLooI0lI<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[23] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && ( (OiOllilOOiI0II0IIilo0IllOOIIIoLii==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OiOllilOOiI0II0IIilo0IllOOIIIoLii<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OLoiILloilO0IIiOOlLoo0LL0ILllliLO>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[24] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && ( (OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[25] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && ( (OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OILlI00OIL0i0OOl0IlOoloII0o0oOlOL>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[26] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && ( (OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OlLIlilLII00OliliLLiLIII0000Ll0o0>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[27] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && ( (OloOLL0I00I0oIIILLo0Ol0Il0lIILL00==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OloOLL0I00I0oIIILLo0Ol0Il0lIILL00<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OooIIILiI0ILoOlO0o0il0LiOoLLLILiO>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[28] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && ( (OioiIOLioLOlOoliOlLli0i0IolIlOLiL==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OioiIOLioLOlOoliOlLli0i0IolIlOLiL<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[29] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && ( (OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OlL0O0LOLillLLIOoOLl0lOOioOiliOol>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[30] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && ( (OiIooILlOili0io0LiiiILIloOi0lIIOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OiIooILlOili0io0LiiiILIloOi0lIIOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OilIIlLl0oo0iilIiiOlilILOlo0IIOOI>=2'd1) ) )) ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[31] <= ( OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && ( (OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) || ( (OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) && (OOI0IILoliiOO0lioiOiO0iloIiOlIlL0>=2'd1) ) )) ;
 OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO <= (OliiILooLoLLIi0IliLO0OO0OOiololoL==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OliiILooLoLLIi0IliLO0OO0OOiololoL<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO>=2'd1) ? 2'd0 : ( OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO+1'd1) ) : OIiol0olIOIoIl0ooOo0OIIi0OOoOLOiO ;
 OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i <= (Oll0lolIi00IiOOiIl00OI0OLoIioOLOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (Oll0lolIi00IiOOiIl00OI0OLoIioOLOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i>=2'd1) ? 2'd0 : ( OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i+1'd1) ) : OIIILoOIoiLL0IoOiLiloOL0ioL0Ll00i ;
 OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo <= (OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo>=2'd1) ? 2'd0 : ( OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo+1'd1) ) : OlLLLLi0i0LlOI00O0IiOOiLI0LL0l0lo ;
 OiLoOlOLii00LILIoloiioLiIoIoioO0L <= (OOOiOlOLli0LLiOOLILIllil0OiLLli0L==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OOOiOlOLli0LLiOOLILIllil0OiLLli0L<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OiLoOlOLii00LILIoloiioLiIoIoioO0L>=2'd1) ? 2'd0 : ( OiLoOlOLii00LILIoloiioLiIoIoioO0L+1'd1) ) : OiLoOlOLii00LILIoloiioLiIoIoioO0L ;
 O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I <= (O0LiLoL0IooiOILoioILLLLli00o0LI0I==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (O0LiLoL0IooiOILoioILLLLli00o0LI0I<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I>=2'd1) ? 2'd0 : ( O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I+1'd1) ) : O00OIO0i0iiIliI0OLoIOLoiIIlIioi0I ;
 OIoLLIoLLLIILi0oi00LolIolIIoliiiI <= (OIolIiLOiOLoO00oiliiollllO0l0OloO==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OIolIiLOiOLoO00oiliiollllO0l0OloO<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OIoLLIoLLLIILi0oi00LolIolIIoliiiI>=2'd1) ? 2'd0 : ( OIoLLIoLLLIILi0oi00LolIolIIoliiiI+1'd1) ) : OIoLLIoLLLIILi0oi00LolIolIIoliiiI ;
 Oi0OollLl0olLol00i0iOOLI0ILliIIIi <= (Oil0OiILooLiiioloiiI0oLLlOlLllo0i==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (Oil0OiILooLiiioloiiI0oLLlOlLllo0i<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((Oi0OollLl0olLol00i0iOOLI0ILliIIIi>=2'd1) ? 2'd0 : ( Oi0OollLl0olLol00i0iOOLI0ILliIIIi+1'd1) ) : Oi0OollLl0olLol00i0iOOLI0ILliIIIi ;
 OO0Ii0IOoilLoILLOIIli0LOLilliLOlI <= (OI0LoL000LIII0lI0LL0LoilIiIlLLiOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OI0LoL000LIII0lI0LL0LoilIiIlLLiOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OO0Ii0IOoilLoILLOIIli0LOLilliLOlI>=2'd1) ? 2'd0 : ( OO0Ii0IOoilLoILLOIIli0LOLilliLOlI+1'd1) ) : OO0Ii0IOoilLoILLOIIli0LOLilliLOlI ;
 O0llOO0ilOIiiioOi0Oloo0IlIILOIlio <= (OoiLi0oolILIllloliLiL0LolIliiLOlo==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OoiLi0oolILIllloliLiL0LolIliiLOlo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((O0llOO0ilOIiiioOi0Oloo0IlIILOIlio>=2'd1) ? 2'd0 : ( O0llOO0ilOIiiioOi0Oloo0IlIILOIlio+1'd1) ) : O0llOO0ilOIiiioOi0Oloo0IlIILOIlio ;
 Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo <= (OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo>=2'd1) ? 2'd0 : ( Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo+1'd1) ) : Oo0LLiO0lOOIl0iIO0lLIiL0ill00OOoo ;
 O0Iliiill00LoolO00Oo0oI00OoolLlLo <= (OioooOOI00ollOl0LiLIl0LIliO00OOii==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OioooOOI00ollOl0LiLIl0LIliO00OOii<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((O0Iliiill00LoolO00Oo0oI00OoolLlLo>=2'd1) ? 2'd0 : ( O0Iliiill00LoolO00Oo0oI00OoolLlLo+1'd1) ) : O0Iliiill00LoolO00Oo0oI00OoolLlLo ;
 O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI <= (OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI>=2'd1) ? 2'd0 : ( O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI+1'd1) ) : O0I0ol0oOLLOLLii0L0IooL0IoiOoLilI ;
 OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O <= (OoolIOILLooLiOLlLiIoO00OooLLL0LLO==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OoolIOILLooLiOLlLiIoO00OooLLL0LLO<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O>=2'd1) ? 2'd0 : ( OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O+1'd1) ) : OOoiOLOioLIlIIOoIo0OOO0Io0OiiIl0O ;
 OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo <= (OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo>=2'd1) ? 2'd0 : ( OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo+1'd1) ) : OliOllLiI0ll0OL0IoIOoLlOOi0lIiLIo ;
 OoILiLOioiOIolLloILoIOLio0iLLoiii <= (OoIIliiLlI0OilooiiILLLOL0oII0ILio==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OoIIliiLlI0OilooiiILLLOL0oII0ILio<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OoILiLOioiOIolLloILoIOLio0iLLoiii>=2'd1) ? 2'd0 : ( OoILiLOioiOIolLloILoIOLio0iLLoiii+1'd1) ) : OoILiLOioiOIolLloILoIOLio0iLLoiii ;
 OLoO0iLi00loILiIo0OlOolilIilOlIii <= (OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OLoO0iLi00loILiIo0OlOolilIilOlIii>=2'd1) ? 2'd0 : ( OLoO0iLi00loILiIo0OlOolilIilOlIii+1'd1) ) : OLoO0iLi00loILiIo0OlOolilIilOlIii ;
 OIIoO0IiLililLIoiilIl00olLoOIlLoL <= (OliilLooOIL0lio0OOioLLoLoLOlioIio==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OliilLooOIL0lio0OOioLLoLoLOlioIio<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OIIoO0IiLililLIoiilIl00olLoOIlLoL>=2'd1) ? 2'd0 : ( OIIoO0IiLililLIoiilIl00olLoOIlLoL+1'd1) ) : OIIoO0IiLililLIoiilIl00olLoOIlLoL ;
 OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo <= (OolioiLoIlIlolO0ooiO0OLOoIlIllIi0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OolioiLoIlIlolO0ooiO0OLOoIlIllIi0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo>=2'd1) ? 2'd0 : ( OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo+1'd1) ) : OiIIOlOlOiI00LI0llIOoo0IOIo00IoOo ;
 OIoI0IOlOLiOllo0iooll00o0lOOoIooo <= (OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OIoI0IOlOLiOllo0iooll00o0lOOoIooo>=2'd1) ? 2'd0 : ( OIoI0IOlOLiOllo0iooll00o0lOOoIooo+1'd1) ) : OIoI0IOlOLiOllo0iooll00o0lOOoIooo ;
 OOLoioilOIOlOOI0iiII0IIOIL0olIL0O <= (OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OOLoioilOIOlOOI0iiII0IIOIL0olIL0O>=2'd1) ? 2'd0 : ( OOLoioilOIOlOOI0iiII0IIOIL0olIL0O+1'd1) ) : OOLoioilOIOlOOI0iiII0IIOIL0olIL0O ;
 OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL <= (O0iiOolLIl0iOLOiLOOLII00IloOo0li0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (O0iiOolLIl0iOLOiLOOLII00IloOo0li0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL>=2'd1) ? 2'd0 : ( OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL+1'd1) ) : OlL0Ooll0lOo0ilLoIOL0lOli0lIIIiIL ;
 OIIi0OoOILoL0LLlLiIOILill0o0ll0OI <= (OLilOOlILoL0oioOOOlOLlOl0li0lIli0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OLilOOlILoL0oioOOOlOLlOl0li0lIli0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OIIi0OoOILoL0LLlLiIOILill0o0ll0OI>=2'd1) ? 2'd0 : ( OIIi0OoOILoL0LLlLiIOILill0o0ll0OI+1'd1) ) : OIIi0OoOILoL0LLlLiIOILill0o0ll0OI ;
 OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo <= (OlIIiOliliiioo0LO0I0IIOIiLLooI0lI==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OlIIiOliliiioo0LO0I0IIOIiLLooI0lI<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo>=2'd1) ? 2'd0 : ( OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo+1'd1) ) : OLLLI0OILilLo0iO0lOo0lO0OlOo00iOo ;
 OLoiILloilO0IIiOOlLoo0LL0ILllliLO <= (OiOllilOOiI0II0IIilo0IllOOIIIoLii==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OiOllilOOiI0II0IIilo0IllOOIIIoLii<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OLoiILloilO0IIiOOlLoo0LL0ILllliLO>=2'd1) ? 2'd0 : ( OLoiILloilO0IIiOOlLoo0LL0ILllliLO+1'd1) ) : OLoiILloilO0IIiOOlLoo0LL0ILllliLO ;
 OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L <= (OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L>=2'd1) ? 2'd0 : ( OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L+1'd1) ) : OOoo0i0LlLlI0LLLo0I0oLoiOio000o0L ;
 OILlI00OIL0i0OOl0IlOoloII0o0oOlOL <= (OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OILlI00OIL0i0OOl0IlOoloII0o0oOlOL>=2'd1) ? 2'd0 : ( OILlI00OIL0i0OOl0IlOoloII0o0oOlOL+1'd1) ) : OILlI00OIL0i0OOl0IlOoloII0o0oOlOL ;
 OlLIlilLII00OliliLLiLIII0000Ll0o0 <= (OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OlLIlilLII00OliliLLiLIII0000Ll0o0>=2'd1) ? 2'd0 : ( OlLIlilLII00OliliLLiLIII0000Ll0o0+1'd1) ) : OlLIlilLII00OliliLLiLIII0000Ll0o0 ;
 OooIIILiI0ILoOlO0o0il0LiOoLLLILiO <= (OloOLL0I00I0oIIILLo0Ol0Il0lIILL00==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OloOLL0I00I0oIIILLo0Ol0Il0lIILL00<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OooIIILiI0ILoOlO0o0il0LiOoLLLILiO>=2'd1) ? 2'd0 : ( OooIIILiI0ILoOlO0o0il0LiOoLLLILiO+1'd1) ) : OooIIILiI0ILoOlO0o0il0LiOoLLLILiO ;
 OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI <= (OioiIOLioLOlOoliOlLli0i0IolIlOLiL==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OioiIOLioLOlOoliOlLli0i0IolIlOLiL<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI>=2'd1) ? 2'd0 : ( OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI+1'd1) ) : OO0ol0lllLOL0OLIlLLOllL0lO0LlOloI ;
 OlL0O0LOLillLLIOoOLl0lOOioOiliOol <= (OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OlL0O0LOLillLLIOoOLl0lOOioOiliOol>=2'd1) ? 2'd0 : ( OlL0O0LOLillLLIOoOLl0lOOioOiliOol+1'd1) ) : OlL0O0LOLillLLIOoOLl0lOOioOiliOol ;
 OilIIlLl0oo0iilIiiOlilILOlo0IIOOI <= (OiIooILlOili0io0LiiiILIloOi0lIIOl==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OiIooILlOili0io0LiiiILIloOi0lIIOl<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OilIIlLl0oo0iilIiiOlilILOlo0IIOOI>=2'd1) ? 2'd0 : ( OilIIlLl0oo0iilIiiOlilILOlo0IIOOI+1'd1) ) : OilIIlLl0oo0iilIiiOlilILOlo0IIOOI ;
 OOI0IILoliiOO0lioiOiO0iloIiOlIlL0 <= (OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00==Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? 2'd0 : (OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00<Oo0olOlL0Oi00o0iLiii0LLOoLIiOilOO) ? ((OOI0IILoliiOO0lioiOiO0iloIiOlIlL0>=2'd1) ? 2'd0 : ( OOI0IILoliiOO0lioiOiO0iloIiOlIlL0+1'd1) ) : OOI0IILoliiOO0lioiOiO0iloIiOlIlL0 ;
 end
 else begin
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 0] <= (OliiILooLoLLIi0IliLO0OO0OOiololoL==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 0] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 1] <= (Oll0lolIi00IiOOiIl00OI0OLoIioOLOl==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 1] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 2] <= (OOoiIiiIiooiO0oLOOIOi0IOOlIiI0o0I==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 2] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 3] <= (OOOiOlOLli0LLiOOLILIllil0OiLLli0L==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 3] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 4] <= (O0LiLoL0IooiOILoioILLLLli00o0LI0I==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 4] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 5] <= (OIolIiLOiOLoO00oiliiollllO0l0OloO==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 5] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 6] <= (Oil0OiILooLiiioloiiI0oLLlOlLllo0i==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 6] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 7] <= (OI0LoL000LIII0lI0LL0LoilIiIlLLiOl==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 7] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 8] <= (OoiLi0oolILIllloliLiL0LolIliiLOlo==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 8] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[ 9] <= (OIOoIiLOIool0iOoO0Ol00i0oiOlllLLO==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[ 9] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[10] <= (OioooOOI00ollOl0LiLIl0LIliO00OOii==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[10] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[11] <= (OIIOllO0iLoIiL0LoLiOlLoILlI00IOOl==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[11] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[12] <= (OoolIOILLooLiOLlLiIoO00OooLLL0LLO==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[12] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[13] <= (OIOLOioO0LLlLl0ioLloiIi0oii0i0lo0==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[13] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[14] <= (OoIIliiLlI0OilooiiILLLOL0oII0ILio==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[14] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[15] <= (OiIOI0LIIiLl0Il0iILOl00IILoiIiO0i==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[15] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[16] <= (OliilLooOIL0lio0OOioLLoLoLOlioIio==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[16] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[17] <= (OolioiLoIlIlolO0ooiO0OLOoIlIllIi0==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[17] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[18] <= (OLiIO0oLOli0Ilo0IlLIolIL0IloilLOo==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[18] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[19] <= (OlIlilOO0L0i0OiI0OlOIOlLlllioLIOo==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[19] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[20] <= (O0iiOolLIl0iOLOiLOOLII00IloOo0li0==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[20] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[21] <= (OLilOOlILoL0oioOOOlOLlOl0li0lIli0==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[21] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[22] <= (OlIIiOliliiioo0LO0I0IIOIiLLooI0lI==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[22] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[23] <= (OiOllilOOiI0II0IIilo0IllOOIIIoLii==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[23] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[24] <= (OOLOOIO0iLOlIIOLoLi0loLi0oIoIOilI==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[24] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[25] <= (OI0LOLOoo00oLLI00LLOLIOlioOLoOl0l==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[25] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[26] <= (OiIOoiLoLlOloIIiLl0l0loL0oloiiIo0==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[26] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[27] <= (OloOLL0I00I0oIIILLo0Ol0Il0lIILL00==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[27] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[28] <= (OioiIOLioLOlOoliOlLli0i0IolIlOLiL==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[28] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[29] <= (OLLoLoiL0lo0IlLolO0lioIiIlIliiLoI==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[29] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[30] <= (OiIooILlOili0io0LiiiILIloOi0lIIOl==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[30] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 O0I0oI0I000LllOOI0L0lOlIl000LIioO[31] <= (OOoLOooiIiLIoiOLO0i0lol0O0Ii0iI00==OO0liOO0iOOIioool0OoLliiiI0l0ilOo)&& OOLIOiLoi0IIOL0LlLliLOILl0ilOIILI[31] && OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 end
 end
 endmodule
 module OlLIiI0ioil0LL0LIOLllLlIiIiOoiL0L ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo , OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI , O0oLi000Lo0oO0oLLoIOllIlo0iOoILio , OiloLLIoolOIiOiOoo00L0I0IOio0lI0L , Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L, OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl, OoIolioOL0iLLOLloI00iIILLiiL0Ooil , OLo0oiiL0ooIliO0I0illLoILiiIoIoOI , OOLOlOo0000iOi0OLOolloLo0iL0iooIi , OLll00OOliOil0O0iLlIooLOLooIIlI0o, OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 , O0li0Illi0oOollo0ooOoIiolOoio0iiL, OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil, OoiloolOiOIoIOolLiOl0OlOiOli0oOOl , OillLliLoolOIiiiILoOILOIloo000iLI , OlLOLoI0iIOLloliOllILlOoIiioOli0L , OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0, OlOiLILOlooo00OLIILLiOioIlO0lLi0l , OiiillOL0OL0oI0O0liIlLIIOL0iLLIli , OlOlO0iLloOIo000llo0LOIloIL0000Li , OIoII0liiOiiO0Lo0illI0iOOI0ll000I , O00iLLLLlOl00oI0loO0OllooooiILolo , /* OiLiiLLIoliLiO0OOloLOlllLiL0ooliI , OilIilioLiOo0Iiioi00OlioIOL0LIOLI , Ol0iIIoo0LoLOIoLiLOOoiil0LoIOiILi , OiI0lioOloloOOIiIOoOLoOOlIl00OI0O , Oil0oLIIoOIOoi0I0iiIIOlL0IiLILOLi , OiIoIlOOioLiILiiIIoLlolllO0ioliLO , OIo0iliLoiiOoLILllILLo0oi0IiiOoLO , Oo0looO00l0oi000oiII00iiiLLL0oOIi , OOLOl0lLLOliOoOlooliOOl0iIL0LOiIL , OI0o0OiiOOioIoIliOIioILoiL0oli0oi , OLillOOlL0II0IiOoOo0lLLILOO00iIoo , OIloLiiOL00oilLo0iiILoOOll0lIlIlO */ OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi, OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 , Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL, OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI );
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo ;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ;
 input O0oLi000Lo0oO0oLLoIOllIlo0iOoILio ;
 input OiloLLIoolOIiOiOoo00L0I0IOio0lI0L ;
 input [3:0] Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L ;
 input [3:0] OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl ;
 input [31:0] OoIolioOL0iLLOLloI00iIILLiiL0Ooil ;
 output [31:0] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi ;
 output [31:0] OLll00OOliOil0O0iLlIooLOLooIIlI0o;
 input [ 15: 0] OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ;
 input [15:0] OoiloolOiOIoIOolLiOl0OlOiOli0oOOl ;
 input [15:0] OillLliLoolOIiiiILoOILOIloo000iLI ;
 input [15:0] OlLOLoI0iIOLloliOllILlOoIiioOli0L ;
 input OlOiLILOlooo00OLIILLiOioIlO0lLi0l ;
 input OiiillOL0OL0oI0O0liIlLIIOL0iLLIli ;
 input OlOlO0iLloOIo000llo0LOIloIL0000Li ;
 input [ 31: 0] OIoII0liiOiiO0Lo0illI0iOOI0ll000I ;
 input [ 1: 0] O00iLLLLlOl00oI0loO0OllooooiILolo ;
 /* input [159: 0] OiLiiLLIoliLiO0OOloLOlllLiL0ooliI ;
 input [ 15: 0] OilIilioLiOo0Iiioi00OlioIOL0LIOLI ;
 output [255: 0] Ol0iIIoo0LoLOIoLiLOOoiil0LoIOiILi ;
 output OiI0lioOloloOOIiIOoOLoOOlIl00OI0O ;
 output Oil0oLIIoOIOoi0I0iiIIOlL0IiLILOLi ;
 output [ 1: 0] OiIoIlOOioLiILiiIIoLlolllO0ioliLO ;
 output OIo0iliLoiiOoLILllILLo0oi0IiiOoLO ;
 input Oo0looO00l0oi000oiII00iiiLLL0oOIi ;
 output OOLOl0lLLOliOoOlooliOOl0iIL0LOiIL ;
 output OI0o0OiiOOioIoIliOIioILoiL0oli0oi ;
 output OLillOOlL0II0IiOoOo0lLLILOO00iIoo ;
 output OIloLiiOL00oilLo0iiILoOOll0lIlIlO ;
 */ output OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi;
 output [255:0] OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 ;
 output Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL;
 input OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI;
 output [63:0] O0li0Illi0oOollo0ooOoIiolOoio0iiL;
 output [31:0] OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil;
 input [31:0] OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0;
 wire [31:0] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 wire [31:0] OO0liOO0iOOIioool0OoLliiiI0l0ilOo;
 wire OiIOLi00lOILlOOL0oLLloL0io0LoIoOL;
 wire [63:0] OoiillIIi0O00lLlIOOiO0OOii0LiLiLO;
 wire [63:0] O0li0Illi0oOollo0ooOoIiolOoio0iiL;
 wire [31:0] OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil;
 wire [15:0] OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ;
 wire [31:0] OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ;
 wire [31:0] OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ;
 wire [31:0] OI00OiLolooiIIiiILoIliO0O0loolIlI ;
 wire [31:0] OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ;
 wire [15:0] OilOOioILlOIIOL0iioIOIi0oloooOoLl ;
 wire OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ;
 wire [ 3: 0] OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ;
 wire OOLOoolOi0LIo0olO0loLllIlllIiiIiI ;
 wire OOOLiLOilooIi0Iio00ilILoLIILOoOoI ;
 wire [ 63: 0] OLLOooI0ILL00ILloiliILLLiioooLliI ;
 wire [ 2: 0] OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ;
 wire [ 15: 0] O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ;
 wire OL0O0IIio0loL0L0Il0li0i00lliIoOOI ;
 wire [4:0] OOLIiil0IlIllLollIl0LIilliOI0iolo;
 wire OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 ;
 wire [3:0] OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI ;
 wire [5:0] OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI ;
 wire OilOOo00lLiOOoiO0ii0oo0oOliOollii ;
 wire [31:0] OIloLiiOL00oilLo0iiILoOOll0lIlIlO ;
 wire [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 wire [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 OOLIoOio0I0i0lliO0OoolLLLLIoLLLlI OO0I0loIlI0iIlIIIOlOLio0oi0lLLLio ( .O0oLi000Lo0oO0oLLoIOllIlo0iOoILio ( O0oLi000Lo0oO0oLLoIOllIlo0iOoILio ) , .OiloLLIoolOIiOiOoo00L0I0IOio0lI0L ( OiloLLIoolOIiOiOoo00L0I0IOio0lI0L ) , .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi), .OlOiLILOlooo00OLIILLiOioIlO0lLi0l ( OlOiLILOlooo00OLIILLiOioIlO0lLi0l ) , .OiiillOL0OL0oI0O0liIlLIIOL0iLLIli ( OiiillOL0OL0oI0O0liIlLIIOL0iLLIli ) , .OL0IIIOOo0000OLoOiO00iiO0lLolLIoO ( OlOlO0iLloOIo000llo0LOIloIL0000Li ) , .OIoII0liiOiiO0Lo0illI0iOOI0ll000I ( OIoII0liiOiiO0Lo0illI0iOOI0ll000I ) , .OlOlLl00OLLOO0ooloIoIli0IIoOLIlOo ( O00iLLLLlOl00oI0loO0OllooooiILolo ) , .OOlOiil0loi0LllL0oOLI00OLoil0l0Ii ( OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ) , .OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI), .O00iLoILoLlOOOolIiiiIOOIlILliLIO0 ( OI00OiLolooiIIiiILoIliO0O0loolIlI ) , .OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl ( OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ) , .OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 ( OilOOioILlOIIOL0iioIOIi0oloooOoLl ) , .OL0Ioll0l0OiIOliOLollLOil000o0iol (OOOLiLOilooIi0Iio00ilILoLIILOoOoI ), .OiILLloIOIIolIio00l00OLOLLIlLoO0o (OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ), .O0LIllilOiLIoilOlLiOio0LiILlllLiI (OOLOoolOi0LIo0olO0loLllIlllIiiIiI ), .OLl0l0oIIoi00000IiiloiLi0OoloLi0L (OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ), .OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO (OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ), .OoOOIil0oLiOILOIIIlIli000O0il000I (OLLOooI0ILL00ILloiliILLLiioooLliI ), .OlLILLOo0IOoilLOO0OlLiioiiioi0IlL (OL0O0IIio0loL0L0Il0li0i00lliIoOOI ), .Olli0loIii0llI00IoOlO0iloLI0oOLOI ( OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ) , .OloOoiioIil00OoLilIliO00IiiillI0I ( O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ) , .OOLIiil0IlIllLollIl0LIilliOI0iolo (OOLIiil0IlIllLollIl0LIilliOI0iolo), .OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI(OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI), .OLOILlOloOoi0OO0oLOOlo0iiIoioilL0(OLOILlOloOoi0OO0oLOOlo0iiIoioilL0), .OLo0oiiL0ooIliO0I0illLoILiiIoIoOI (OLo0oiiL0ooIliO0I0illLoILiiIoIoOI), .OO0liOO0iOOIioool0OoLliiiI0l0ilOo (OO0liOO0iOOIioool0OoLliiiI0l0ilOo), .OiIOLi00lOILlOOL0oLLloL0io0LoIoOL (OiIOLi00lOILlOOL0oLLloL0io0LoIoOL), .OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI(OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI) , .OilOOo00lLiOOoiO0ii0oo0oOliOollii (OilOOo00lLiOOoiO0ii0oo0oOliOollii) , .OIloLiiOL00oilLo0iiILoOOll0lIlIlO ( OIloLiiOL00oilLo0iiILoOOll0lIlIlO ) , .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl), .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol), .OoiillIIi0O00lLlIOOiO0OOii0LiLiLO (OoiillIIi0O00lLlIOOiO0OOii0LiLiLO), .OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil (OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil), .OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0 (OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0), .OLll00OOliOil0O0iLlIooLOLooIIlI0o(OLll00OOliOil0O0iLlIooLOLooIIlI0o), .O0li0Illi0oOollo0ooOoIiolOoio0iiL (O0li0Illi0oOollo0ooOoIiolOoio0iiL) );
 OILLilL0iiliiLLO0IL0LiOoLILlOL0iO OILLilL0iiliiLLO0IL0LiOoLILlOL0iO ( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo ) , .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ( OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI ) , .Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L (Ooo00loiOoLioL0O0LoOlLio0oI0lIo0L), .OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl (OII00ILLo0I0I0lLlo0LLi0o0i0L0LIOl), .OoIolioOL0iLLOLloI00iIILLiiL0Ooil (OoIolioOL0iLLOLloI00iIILLiiL0Ooil), .OOLIiil0IlIllLollIl0LIilliOI0iolo (OOLIiil0IlIllLollIl0LIilliOI0iolo), .OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI(OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI), .OLOILlOloOoi0OO0oLOOlo0iiIoioilL0(OLOILlOloOoi0OO0oLOOlo0iiIoioilL0), .OLll00OOliOil0O0iLlIooLOLooIIlI0o(OLll00OOliOil0O0iLlIooLOLooIIlI0o), .OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI(OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI) , .OilOOo00lLiOOoiO0ii0oo0oOliOollii (OilOOo00lLiOOoiO0ii0oo0oOliOollii) , .OolIOLOooiLLIllI0LOLIolllLoilolIl (OolIOLOooiLLIllI0LOLIolllLoilolIl), .O0IOooLliOlIllOliILoolIIoIiO0Ilol (O0IOooLliOlIllOliILoolIIoIiO0Ilol), .OLo0oiiL0ooIliO0I0illLoILiiIoIoOI (OLo0oiiL0ooIliO0I0illLoILiiIoIoOI), .OO0liOO0iOOIioool0OoLliiiI0l0ilOo (OO0liOO0iOOIioool0OoLliiiI0l0ilOo), .OiIOLi00lOILlOOL0oLLloL0io0LoIoOL (OiIOLi00lOILlOOL0oLLloL0io0LoIoOL), .OOLOlOo0000iOi0OLOolloLo0iL0iooIi (OOLOlOo0000iOi0OLOolloLo0iL0iooIi), .OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 (OL0lOiIIlLoILOLIIiIoLoLOILl0LOO00 ) , .OoiloolOiOIoIOolLiOl0OlOiOli0oOOl (OoiloolOiOIoIOolLiOl0OlOiOli0oOOl), .OillLliLoolOIiiiILoOILOIloo000iLI (OillLliLoolOIiiiILoOILOIloo000iLI), .OlLOLoI0iIOLloliOllILlOoIiioOli0L (OlLOLoI0iIOLloliOllILlOoIiioOli0L), .OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ( OliIO0oOoLIi0il0LLooL0Oo00Lo0lOoI ) , .OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ( OoiOoloi0I0IL00Ii0LIO0LOLIllIOIII ) , .OOLOoolOi0LIo0olO0loLllIlllIiiIiI ( OOLOoolOi0LIo0olO0loLllIlllIiiIiI ) , .OOOLiLOilooIi0Iio00ilILoLIILOoOoI ( OOOLiLOilooIi0Iio00ilILoLIILOoOoI ) , .OLLOooI0ILL00ILloiliILLLiioooLliI ( OLLOooI0ILL00ILloiliILLLiioooLliI ) , .OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ( OILoli0OIOIIOI0OiliOo0i0OLoliOOiI ) , .O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ( O0olOiI0OOI0OOIOOiI0L0OiLLLOo0OlI ) , .OL0O0IIio0loL0L0Il0li0i00lliIoOOI ( OL0O0IIio0loL0L0Il0li0i00lliIoOOI ) , .OilOOioILlOIIOL0iioIOIi0oloooOoLl ( OilOOioILlOIIOL0iioIOIi0oloooOoLl ) , .OI00OiLolooiIIiiILoIliO0O0loolIlI ( OI00OiLolooiIIiiILoIliO0O0loolIlI ) , .OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ( OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo ) , .OIloLiiOL00oilLo0iiILoOOll0lIlIlO ( OIloLiiOL00oilLo0iiILoOOll0lIlIlO ) , .OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ( OOLOIoLliliO0Li0OLlIO0OOL0Ollio0O ) , .OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI ( OIlLi0iolo0LIOI0o00OooIOOL0O0oOLI), .OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ( OIIOLLOIlOlLoi0oiOioLilOiioiiliLO ) , .OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi (OOiLOIIllLlOO0iLIiLol0IIOOLIOiOOi), .OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 (OLOILliLL0OlLIo0ol0IIlliOLiL0i0O0 ), .Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL (Oo0ILIoiL0oI0OOo0OL0ioIiOlLoiiOIL), .OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI (OOIllIlIIIO0LOOo0LoOilloIoIIOLOLI) );
 endmodule
 module OoILi0OOLIloI0O0lO0lOLo0iLlO0o0oo ( Ol00oIollLiioLLLoiOiolOL00iiOlIoo, OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI, OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL, OO0o0l0ioiI0oo0oiOL00LooiIIoli00o, OollLiiii0o0lIiIiL0OL0OLiLllLL0I0, OoIlOoIlIooO0lIIooIoillLl0O0OLlol, OOLOOIi000oLlOiO0LLiIIIoIIO0ILool, OOlOiil0loi0LllL0oOLI00OLoil0l0Ii, OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl, Olli0loIii0llI00IoOlO0iloLI0oOLOI, OloOoiioIil00OoLilIliO00IiiillI0I, O00iLoILoLlOOOolIiiiIOOIlILliLIO0, OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl, OL0Ioll0l0OiIOliOLollLOil000o0iol, OoOOIil0oLiOILOIIIlIli000O0il000I, OiILLloIOIIolIio00l00OLOLLIlLoO0o, OLl0l0oIIoi00000IiiloiLi0OoloLi0L, O0LIllilOiLIoilOlLiOio0LiILlllLiI, OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO, OiIoiiOIOOi0OLILo0oIOOioO0IioLI00, OiLIiLoILI0LiLOlLIoOolOolIIlOIllI, OiiiIllliL0oLoOIliliIilLiollooiII , OI0ioooOlLlIoLiL0IO0oOII0OlLiOo0I , O0lOOlIOlIo0IILillLi0liOLlO00OILL , OILLO0olLiLlOoOolOloOOLiliIIiIOLO , OIiOoioOIOoLIOO0OLioll0I0IIiIoOOi , OOIOlI0OolOlLlOOIii0ioo00iio0IIil , OIloLiiOL00oilLo0iiILoOOll0lIlIlO , OLo0oiiL0ooIliO0I0illLoILiiIoIoOI , OO0liOO0iOOIioool0OoLliiiI0l0ilOo , OiIOLi00lOILlOOL0oLLloL0io0LoIoOL , OoiillIIi0O00lLlIOOiO0OOii0LiLiLO, OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil, OLll00OOliOil0O0iLlIooLOLooIIlI0o, OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0, O0li0Illi0oOollo0ooOoIiolOoio0iiL );
 localparam [2:0] IDLE = 3'b000;
 localparam [2:0] PARSE = 3'b001;
 localparam [2:0] PAYLOAD_OUT = 3'b011;
 localparam [2:0] SEARCH = 3'b010;
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI;
 input OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL;
 input [63:0] OO0o0l0ioiI0oo0oiOL00LooiIIoli00o;
 input OollLiiii0o0lIiIiL0OL0OLiLllLL0I0;
 input OoIlOoIlIooO0lIIooIoillLl0O0OLlol;
 input [2:0] OOLOOIi000oLlOiO0LLiIIIoIIO0ILool;
 input [31:0] OOlOiil0loi0LllL0oOLI00OLoil0l0Ii;
 input [31:0] OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl;
 output [15:0] Olli0loIii0llI00IoOlO0iloLI0oOLOI;
 output [15:0] OloOoiioIil00OoLilIliO00IiiillI0I;
 output [31:0] O00iLoILoLlOOOolIiiiIOOIlILliLIO0;
 output [31:0] OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl;
 output OL0Ioll0l0OiIOliOLollLOil000o0iol;
 output [63:0] OoOOIil0oLiOILOIIIlIli000O0il000I;
 output OiILLloIOIIolIio00l00OLOLLIlLoO0o;
 output [3:0] OLl0l0oIIoi00000IiiloiLi0OoloLi0L;
 output O0LIllilOiLIoilOlLiOio0LiILlllLiI;
 output [2:0] OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO;
 output [15:0] OiIoiiOIOOi0OLILo0oIOOioO0IioLI00;
 input [4:0] OiLIiLoILI0LiLOlLIoOolOolIIlOIllI;
 input OiiiIllliL0oLoOIliliIilLiollooiII ;
 input [3:0] OI0ioooOlLlIoLiL0IO0oOII0OlLiOo0I ;
 input [15:0] O0lOOlIOlIo0IILillLi0liOLlO00OILL ;
 input [ 5:0] OILLO0olLiLlOoOolOloOOLiliIIiIOLO ;
 input [5:0] OIiOoioOIOoLIOO0OLioll0I0IIiIoOOi ;
 input OOIOlI0OolOlLlOOIii0ioo00iio0IIil ;
 input [31:0] OIloLiiOL00oilLo0iiILoOOll0lIlIlO ;
 input [31:0 ] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 input [31:0 ] OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 input OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 output [63:0] OoiillIIi0O00lLlIOOiO0OOii0LiLiLO;
 output [31:0] OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil;
 input [31:0] OLll00OOliOil0O0iLlIooLOLooIIlI0o;
 input [31:0] OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0;
 output [63:0] O0li0Illi0oOollo0ooOoIiolOoio0iiL;
 reg [63:0] OoiillIIi0O00lLlIOOiO0OOii0LiLiLO;
 reg [31:0] OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil;
 reg [63:0] O0li0Illi0oOollo0ooOoIiolOoio0iiL;
 reg [15:0] OloOoiioIil00OoLilIliO00IiiillI0I;
 reg [31:0] O00iLoILoLlOOOolIiiiIOOIlILliLIO0;
 reg [31:0] OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl;
 reg OL0Ioll0l0OiIOliOLollLOil000o0iol;
 reg [63:0] OoOOIil0oLiOILOIIIlIli000O0il000I;
 reg OiILLloIOIIolIio00l00OLOLLIlLoO0o;
 reg [3:0] OLl0l0oIIoi00000IiiloiLi0OoloLi0L;
 reg O0LIllilOiLIoilOlLiOio0LiILlllLiI;
 reg [2:0] OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO;
 reg [15:0] OiIoiiOIOOi0OLILo0oIOOioO0IioLI00;
 reg [2:0] Olo0I0OOli0Oii0IoOOLloiiliollIolO;
 reg [2:0] OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL;
 reg [103:0] fivetuple_pre [0:31] ;
 reg [103:0] OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli = 104'b0;
 reg [135:0] fivetuple_seq_pre [0:31] ;
 wire [135:0] OlIIIll00io0lOLOioI0IOilLLoOIoO0l ;
 reg [135:0] OO0iOiIoo0OLLILiLolOIOoIlIIolIOoL;
 reg [31:0] OLlOOLliiiLol0illoioo0LOoOOllo0O0 = {32{1'b0}};
 reg [31:0] OI00llolIOiOLO0I0OioOOIlilLi0lILi = {32{1'b0}};
 wire [31:0] Oi0iol0looOo0iLo0LIiOLloiIloOoOol;
 wire [31:0] OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo;
 reg OOioolL0l0iLOiO00iiIlIiOIOOOL000L;
 reg O00ioIooO0looL0lL0lil0ooIIOliIl0L;
 reg OOo0loo0OOILILoOl0LoiLOi0ILIoOOLO;
 wire OIiiO0OILoiioIoILoLoIioooOolOOioL;
 reg O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll;
 reg OIl0iO0LoI0olLLoIoLiloOiLLliLiLol = 1'd0 ;
 reg OIOLLioLILi0o0iiLIo0IOLIOoO0liioi = 1'd0 ;
 reg OlOliIi0llill0LolIOiLoLloLIllIlIO;
 reg [31:0] OLOiOL0L0LOiloiIIOliIOioioIOOLOOi;
 reg [31:0] Ol0LLOl0OOlilLOiiLLill0OIlLil0iLI;
 reg [7:0] O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0;
 reg [15:0] OIllLolLlliOllI00ioL0LloL0OiLIIIL;
 reg [15:0] OLLLoLiIIlILoOloIilLO0oIlOloOILOO;
 reg OoiIoiOllllIL0OOIOO0OlLIOIIolIloi;
 wire [15:0] OoOIIlLLOIOIiloOi0oO0OliLllILoOIo;
 reg [15:0] OL0I0LLIIli0LOLliOIol00OLioi0l0Li;
 reg [5:0] OiOiioOOIOLL0OO000O0iLiiLILLII0ii;
 reg [5:0] OO0OIooOL0O0o0O0lL0OO0oOiiOIO00Io;
 reg [6:0] OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi;
 reg O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI;
 reg [6:0] OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo;
 reg O0L00liiLLLiiL00OlOoOilOOiil00LIl;
 reg OLiLiILlL0IOoloIIlooioOLIiOOoOloi;
 reg [31:0] OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo;
 reg [31:0] O0iO0LoL0OllIoILOLLlioliIiIoOIl0i;
 wire [31:0] OLLi0iLioIOLL0LL0lIL0lIIlL0LI0l0L;
 reg [5:0] O0iILILLiIlLLIOlOolIL0LOiLlIio0Ii;
 reg OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 ;
 reg Oli0IIIlllIiO0llio0OOLliOIiOLiioL;
 reg [63:0] OiOIIO0ol0IOIoLIO0ililo0lloOlIiII;
 reg [63:0] OLiOLOo0IiliIiiIlil0olIlIlooi0IoL;
 reg O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo;
 reg [63:0] OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0;
 reg [63:0] OoLILillIiOiooIoIoLLilL0Llooi0OlI;
 wire OlOiLILOlooo00OLIILLiOioIlO0lLi0l;
 wire OiiillOL0OL0oI0O0liIlLIIOL0iLLIli;
 reg [15:0] OiiiiiOOI0lloLLIILlOOlolLlLo0olLL;
 reg OLOIl0loioiIllIlOlOLiOO0ooiiLliio;
 reg [2:0] OIIILilLlLLiolIILLOilOllLili00LoI;
 reg [11:0] OIOll0OLlLIloLlIOiLi0lo0olOIoOOII = 12'd0;
 assign OlOiLILOlooo00OLIILLiOioIlO0lLi0l = OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL & OollLiiii0o0lIiIiL0OL0OLiLllLL0I0;
 assign OiiillOL0OL0oI0O0liIlLIIOL0iLLIli = OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL & OoIlOoIlIooO0lIIooIoillLl0O0OLlol;
 always @ (posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0 <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o;
 OoLILillIiOiooIoIoLLilL0Llooi0OlI <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0;
 end
 always @ (posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OIOll0OLlLIloLlIOiLi0lo0olOIoOOII <= 12'd0;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OIOll0OLlLIloLlIOiLi0lo0olOIoOOII <= OIOll0OLlLIloLlIOiLi0lo0olOIoOOII + 12'd8;
 reg [15:0] OIIOLLOIlOlLoi0oiOioLilOiioiiliLO;
 assign Olli0loIii0llI00IoOlO0iloLI0oOLOI = OL0I0LLIIli0LOLliOIol00OLioi0l0Li - OiOiioOOIOLL0OO000O0iLiiLILLII0ii - OO0OIooOL0O0o0O0lL0OO0oOiiOIO00Io;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) Olo0I0OOli0Oii0IoOOLloiiliollIolO <= IDLE;
 else Olo0I0OOli0Oii0IoOOLloiiliollIolO <= OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL;
 always @(*) case(Olo0I0OOli0Oii0IoOOLloiiliollIolO) IDLE: begin
 if(OlOiLILOlooo00OLIILLiOioIlO0lLi0l) OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = PARSE;
 else OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = IDLE;
 end
 PARSE: begin
 if(!OIl0iO0LoI0olLLoIoLiloOiLLliLiLol || !OIOLLioLILi0o0iiLIo0IOLIOoO0liioi ) OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = IDLE;
 else if(OoiIoiOllllIL0OOIOO0OlLIOIIolIloi&&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 if(|Oi0iol0looOo0iLo0LIiOLloiIloOoOol) OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = PAYLOAD_OUT;
 else OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = SEARCH;
 end
 else OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = PARSE;
 end
 PAYLOAD_OUT: begin
 if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = IDLE;
 else OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = PAYLOAD_OUT;
 end
 SEARCH: begin
 if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = IDLE;
 else OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = SEARCH;
 end
 default: OlIIIilOLiLlIOoLi0iLo0oLLOiIiilLL = IDLE;
 endcase generate genvar ch;
 for(ch = 0;
 ch < 32;
 ch=ch+1) begin
: O0IliOLIlIOLlOIoioi0OlIL0IOliiIol always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if((fivetuple_seq_pre[ch] == OlIIIll00io0lOLOioI0IOilLLoOIoO0l)&& OI00llolIOiOLO0I0OioOOIlilLi0lILi[ch]&&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OLlOOLliiiLol0illoioo0LOoOOllo0O0[ch] <= 1'b0;
 else if (OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl[ch]) OLlOOLliiiLol0illoioo0LOoOOllo0O0[ch] <= 1'b0;
 else if(OOlOiil0loi0LllL0oOLI00OLoil0l0Ii[ch]) OLlOOLliiiLol0illoioo0LOoOOllo0O0[ch] <= 1'b1;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OOlOiil0loi0LllL0oOLI00OLoil0l0Ii[ch]) fivetuple_seq_pre[ch] <= OO0iOiIoo0OLLILiLolOIOoIlIIolIOoL;
 end
 assign Oi0iol0looOo0iLo0LIiOLloiIloOoOol[ch] = OLlOOLliiiLol0illoioo0LOoOOllo0O0[ch] && (fivetuple_seq_pre[ch] == OlIIIll00io0lOLOioI0IOilLLoOIoO0l) && OI00llolIOiOLO0I0OioOOIlilLi0lILi[ch]&&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL;
 assign OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo[ch] = OLlOOLliiiLol0illoioo0LOoOOllo0O0[ch] && (fivetuple_seq_pre[ch][103:0] == OlIIIll00io0lOLOioI0IOilLLoOIoO0l[103:0])&&(fivetuple_seq_pre[ch][135:104] != OlIIIll00io0lOLOioI0IOilLLoOIoO0l[135:104]) && OI00llolIOiOLO0I0OioOOIlilLi0lILi[ch]&& OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) O00iLoILoLlOOOolIiiiIOOIlILliLIO0[ch] <= 1'b0;
 else if(O0LIllilOiLIoilOlLiOio0LiILlllLiI&&OL0Ioll0l0OiIOliOLollLOil000o0iol) O00iLoILoLlOOOolIiiiIOOIlILliLIO0[ch] <= 1'b0;
 else if(Oi0iol0looOo0iLo0LIiOLloiIloOoOol[ch]) O00iLoILoLlOOOolIiiiIOOIlILliLIO0[ch] <= 1'b1;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl[ch] <= 1'b0;
 else if(O0LIllilOiLIoilOlLiOio0LiILlllLiI&&OL0Ioll0l0OiIOliOLollLOil000o0iol) OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl[ch] <= 1'b0;
 else if(OL0O0oOlll0oOoLiioOiLl00oiIlLOoIo[ch]) OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl[ch] <= 1'b1;
 end
 end
 endgenerate reg [7:0] OillLLIloOooLolooI0oiLLOO0LOoliio = 8'b0;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OillLLIloOooLolooI0oiLLOO0LOoliio <= 8'b0;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OillLLIloOooLolooI0oiLLOO0LOoliio <= OillLLIloOooLolooI0oiLLOO0LOoliio + 1'b1;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd1)) begin
 if(OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[31:16]==16'h8100) O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll <= 1'b1;
 else O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll <= 1'b0;
 end
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OOioolL0l0iLOiO00iiIlIiOIOOOL000L <= 1'b0;
 else if(O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll && OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd2)&& (OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]== 16'h0800)) OOioolL0l0iLOiO00iiIlIiOIOOOL000L <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd1) && (OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[31:16]== 16'h0800)) OOioolL0l0iLOiO00iiIlIiOIOOOL000L <= 1'b1;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3)) begin
 if(!OOioolL0l0iLOiO00iiIlIiOIOOOL000L) OIl0iO0LoI0olLLoIoLiloOiLLliLiLol <= 1'b0;
 else OIl0iO0LoI0olLLoIoLiloOiLLliLiLol <= 1'b1;
 end
 else OIl0iO0LoI0olLLoIoLiloOiLLliLiLol <= 1'b1;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) O00ioIooO0looL0lL0lil0ooIIOliIl0L <= 1'b0;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd2)&&(OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[7:0]== 8'h06)) O00ioIooO0looL0lL0lil0ooIIOliIl0L <= 1'b1;
 end
 reg OiIlilLLlL0IIL0OoLLoOOoLoiLo0LiIO;
 always @(*) begin
 if(O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll && OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3)&&(OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[39:32]== 8'h06)) OiIlilLLlL0IIL0OoLLoOOoLoiLo0LiIO = 1'b1;
 else OiIlilLLlL0IIL0OoLLoOOoLoiLo0LiIO = 1'b0;
 end
 always @ (posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OOo0loo0OOILILoOl0LoiLOi0ILIoOOLO <= 1'b0;
 else if(OiIlilLLlL0IIL0OoLLoOOoLoiLo0LiIO) OOo0loo0OOILILoOl0LoiLOi0ILIoOOLO <= 1'b1;
 assign OIiiO0OILoiioIoILoLoIioooOolOOioL = OOo0loo0OOILILoOl0LoiLOi0ILIoOOLO | OiIlilLLlL0IIL0OoLLoOOoLoiLo0LiIO | O00ioIooO0looL0lL0lil0ooIIOliIl0L;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3)) begin
 if(!OIiiO0OILoiioIoILoLoIioooOolOOioL) OIOLLioLILi0o0iiLIo0IOLIOoO0liioi <= 1'b0;
 else OIOLLioLILi0o0iiLIo0IOLIOoO0liioi <= 1'b1;
 end
 else begin
 OIOLLioLILi0o0iiLIo0IOLIOoO0liioi <= 1'b1;
 end
 end
 wire OliO0illloo0lOoOOioOiO0lIlOLL0ILI;
 assign OliO0illloo0lOoOOioOiO0lIlOLL0ILI = OOioolL0l0iLOiO00iiIlIiOIOOOL000L && !O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd1) && (OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[31:16]== 16'h0800))begin
 OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[11:8],2'b00} + 7'd14;
 OiOiioOOIOLL0OO000O0iLiiLILLII0ii <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[11:8],2'b00};
 end
 else if(O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll && OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd2) && (OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]== 16'h0800)) begin
 OiOiioOOIOLL0OO000O0iLiiLILLII0ii <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[43:40],2'b00};
 OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[43:40],2'b00} + 7'd18;
 end
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OliO0illloo0lOoOOioOiO0lIlOLL0ILI) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd2) begin
 O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0 <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[7:0];
 OL0I0LLIIli0LOLliOIol00OLioi0l0Li <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48];
 end
 else if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3) begin
 OLOiOL0L0LOiloiIIOliIOioioIOOLOOi <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16];
 end
 else if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd4) begin
 Ol0LLOl0OOlilLOiiLLill0OIlLil0iLI <= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 end
 end
 else if(O0o0Lo00oOl0LL0lLiOI00I00i0oLo0Ll) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd2) begin
 OL0I0LLIIli0LOLliOIol00OLioi0l0Li <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[31:16];
 end
 else if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3) begin
 O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0 <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[39:32];
 end
 else if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd4) begin
 Ol0LLOl0OOlilLOiiLLill0OIlLil0iLI <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16];
 OLOiOL0L0LOiloiIIOliIOioioIOOLOOi <= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 end
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 if ( ~OIiiO0OILoiioIoILoLoIioooOolOOioL || ~OOioolL0l0iLOiO00iiIlIiOIOOOL000L ) begin
 O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'd0 ;
 end
 else begin
 case(OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi[6:3]) 4'd4: begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 4'd5: begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd4)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 4'd6: begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd5)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 4'd7: begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd6)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 4'd8: begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd7)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 4'd9: begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd8)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 default : begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd3)) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b1;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI <= 1'b0;
 end
 endcase end
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) begin
 OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 <= 1'b0;
 Oli0IIIlllIiO0llio0OOLliOIiOLiioL <= 1'b0;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 <= O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI ;
 Oli0IIIlllIiO0llio0OOLliOIiOLiioL <= OOLLO0Oii00IOO0OloOoolIOiLLilIiI0;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) case(OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi[2:0]) 3'b010: begin
 if(O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 if(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd4) OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli <= {OLOiOL0L0LOiloiIIOliIOioioIOOLOOi,OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48],O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0,OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16]};
 else OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli <= {OLOiOL0L0LOiloiIIOliIOioioIOOLOOi,Ol0LLOl0OOlilLOiiLLill0OIlLil0iLI,O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0,OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16]};
 end
 end
 3'b110: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli <= {OLOiOL0L0LOiloiIIOliIOioioIOOLOOi,Ol0LLOl0OOlilLOiiLLill0OIlLil0iLI,O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0,OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 end
 default: begin
 if(O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli <= {OLOiOL0L0LOiloiIIOliIOioioIOOLOOi,Ol0LLOl0OOlilLOiiLLill0OIlLil0iLI,O0oOLOOOiOL0LIiolIoIlOLlOoOlLLOl0,OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16]};
 end
 end
 endcase always @(*) case(OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi[2:0]) 3'b010: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo = {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 else begin
 OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo = 32'd0;
 end
 end
 3'b110: begin
 if(Oli0IIIlllIiO0llio0OOLliOIiOLiioL & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[47:16]};
 end
 else begin
 OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo = 32'd0;
 end
 end
 default: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo = {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 else begin
 OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo = 32'd0;
 end
 end
 endcase assign OLLi0iLioIOLL0LL0lIL0lIIlL0LI0l0L = O0iO0LoL0OllIoILOLLlioliIiIoOIl0i + Olli0loIii0llI00IoOlO0iloLI0oOLOI;
 assign OlIIIll00io0lOLOioI0IOilLLoOIoO0l = {OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli,OLIOoOIiOoliLl0IOiLIiiolilIiOIoOo};
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) OO0iOiIoo0OLLILiLolOIOoIlIIolIOoL <= {OoiLIlLoIiOlL0OOl0LOLill0Il0OLOli,OLLi0iLioIOLL0LL0lIL0lIIlL0LI0l0L};
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OoiIoiOllllIL0OOIOO0OlLIOIIolIloi <= 1'b0;
 else begin
 case(OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi[2:0]) 3'b010: begin
 if(O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OoiIoiOllllIL0OOIOO0OlLIOIIolIloi <= 1'b1;
 end
 end
 3'b110: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0&&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OoiIoiOllllIL0OOIOO0OlLIOIIolIloi <= 1'b1;
 end
 end
 default: begin
 if(O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OoiIoiOllllIL0OOIOO0OlLIOIIolIloi <= 1'b1;
 end
 end
 endcase end
 reg [6:0] O0Ll0IiOilIO0iiLiiiliLoILL0ILiLlo;
 always @ (posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 O0Ll0IiOilIO0iiLiiiliLoILL0ILiLlo <= OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi;
 end
 generate genvar chn;
 for(chn = 0;
 chn < 32;
 chn=chn+1) begin
: OIIi0oo0l0OOI00iIlOl0oiOLoLi0OoLi always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OOlOiil0loi0LllL0oOLI00OLoil0l0Ii[chn] && !O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI) OI00llolIOiOLO0I0OioOOIlilLi0lILi[chn] <= 1'b0;
 else if(OLlOOLliiiLol0illoioo0LOoOOllo0O0[chn] | OOlOiil0loi0LllL0oOLI00OLoil0l0Ii[chn]) begin
 case(OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi[2:0]) 3'b010: begin
 if(O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OI00llolIOiOLO0I0OioOOIlilLi0lILi[chn] <= 1'b1;
 end
 end
 3'b110: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0&&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OI00llolIOiOLO0I0OioOOIlilLi0lILi[chn] <= 1'b1;
 end
 end
 default: begin
 if(O0ioIL0IOLLlOoLiIOolLIlLo0ioIILiI & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL ) begin
 OI00llolIOiOLO0I0OioOOIlilLi0lILi[chn] <= 1'b1;
 end
 end
 endcase end
 else OI00llolIOiOLO0I0OioOOIlilLi0lILi[chn] <= 1'b0;
 end
 endgenerate always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) begin
 OLiLiILlL0IOoloIIlooioOLIiOOoOloi <= 1'b0;
 end
 else begin
 case(OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi[2:0]) 3'b010: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OIllLolLlliOllI00ioL0LloL0OiLIIIL <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[47:32];
 OLLLoLiIIlILoOloIilLO0oIlOloOILOO <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[31:16];
 OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[15:12],2'b00} + OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi;
 OLiLiILlL0IOoloIIlooioOLIiOOoOloi <= 1'b1;
 OO0OIooOL0O0o0O0lL0OO0oOiiOIO00Io <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[15:12],2'b00};
 O0iO0LoL0OllIoILOLLlioliIiIoOIl0i <= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 end
 3'b110: begin
 if(Oli0IIIlllIiO0llio0OOLliOIiOLiioL & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) begin
 OIllLolLlliOllI00ioL0LloL0OiLIIIL <= OoLILillIiOiooIoIoLLilL0Llooi0OlI[15:0];
 OLLLoLiIIlILoOloIilLO0oIlOloOILOO <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[63:48];
 OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:44],2'b00} + OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi;
 OLiLiILlL0IOoloIIlooioOLIiOOoOloi <= 1'b1;
 OO0OIooOL0O0o0O0lL0OO0oOiiOIO00Io <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:44],2'b00};
 O0iO0LoL0OllIoILOLLlioliIiIoOIl0i <= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[47:16]};
 end
 end
 default: begin
 if(OOLLO0Oii00IOO0OloOoolIOiLLilIiI0 & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL ) begin
 OIllLolLlliOllI00ioL0LloL0OiLIIIL <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[47:32];
 OLLLoLiIIlILoOloIilLO0oIlOloOILOO <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[31:16];
 OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[15:12],2'b00} + OIiLLI0OOO0loOl0lII0i0oIiLOOIlLoi;
 OLiLiILlL0IOoloIIlooioOLIiOOoOloi <= 1'b1;
 OO0OIooOL0O0o0O0lL0OO0oOiiOIO00Io <= {OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[15:12],2'b00};
 O0iO0LoL0OllIoILOLLlioliIiIoOIl0i <= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]};
 end
 end
 endcase end
 always @(*) begin
 case(OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo[6:3]) 4'd6: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi && OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd6)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd7: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd7)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd8: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd8)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd9: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd9)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd10: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd10)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd11: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd11)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd4: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd4)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd5: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd5)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd12: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd12)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 4'd13: begin
 if(OLiLiILlL0IOoloIIlooioOLIiOOoOloi &&OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd13)) O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b1;
 else O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 default : begin
 O0L00liiLLLiiL00OlOoOilOOiil00LIl = 1'b0;
 end
 endcase end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli & O0L00liiLLLiiL00OlOoOilOOiil00LIl & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OloOoiioIil00OoLilIliO00IiiillI0I <= 4'd8 - OOLOOIi000oLlOiO0LLiIIIoIIO0ILool - OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo[2:0];
 else if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OloOoiioIil00OoLilIliO00IiiillI0I <= OloOoiioIil00OoLilIliO00IiiillI0I + (4'd8 - OOLOOIi000oLlOiO0LLiIIIoIIO0ILool);
 else if(O0L00liiLLLiiL00OlOoOilOOiil00LIl & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OloOoiioIil00OoLilIliO00IiiillI0I <= 4'd8 - OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo[2:0];
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OloOoiioIil00OoLilIliO00IiiillI0I <= OloOoiioIil00OoLilIliO00IiiillI0I + 4'd8;
 always @(*) if(Olo0I0OOli0Oii0IoOOLloiiliollIolO == SEARCH) begin
 if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[47:32],OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd2;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[39:24],OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[7:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:40]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd3;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[31:16],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:32]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd4;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[23:8],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[55:24]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd5;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd6;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[7:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:56],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[39:8]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd7;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[63:48],OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[31:0]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd0;
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[55:40],OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[23:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:56]}== 48'h02000100044c)) begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b1;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd1;
 end
 else begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b0;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd0;
 end
 end
 else begin
 OLOIl0loioiIllIlOlOLiOO0ooiiLliio = 1'b0;
 OIIILilLlLLiolIILLOilOllLili00LoI = 3'd0;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[31:16];
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[7:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:40]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[23:8];
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:32]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[15:0];
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[55:24]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= {OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[7:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:56]};
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[47:16]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:48];
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[39:8]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[55:40];
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[31:0]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[47:32];
 end
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && ({OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[23:0],OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[63:56]}== 32'h0100044c)) begin
 OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 <= OLlI0OL0ILioILoOLOOOOLoOooIOLl0L0[39:24];
 end
 reg OLi00LI00i0LIIiO0olIo00Liii0ILLii = 1'b0;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(Olo0I0OOli0Oii0IoOOLloiiliollIolO == PAYLOAD_OUT) begin
 OiILLloIOIIolIio00l00OLOLLIlLoO0o <= O0L00liiLLLiiL00OlOoOilOOiil00LIl;
 OLl0l0oIIoi00000IiiloiLi0OoloLi0L <= OLiO0OLOlLI0OIlOlilLiiOloOOiOLiLo[2:0];
 OL0Ioll0l0OiIOliOLollLOil000o0iol <= OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL & (O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo|O0L00liiLLLiiL00OlOoOilOOiil00LIl);
 OoOOIil0oLiOILOIIIlIli000O0il000I <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o;
 end
 else if(Olo0I0OOli0Oii0IoOOLloiiliollIolO == SEARCH) begin
 OiILLloIOIIolIio00l00OLOLLIlLoO0o <= OLOIl0loioiIllIlOlOLiOO0ooiiLliio & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL && (OLi00LI00i0LIIiO0olIo00Liii0ILLii == 1'b0);
 OLl0l0oIIoi00000IiiloiLi0OoloLi0L <= OIIILilLlLLiolIILLOilOllLili00LoI;
 OL0Ioll0l0OiIOliOLollLOil000o0iol <= OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL & (O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo | OLOIl0loioiIllIlOlOLiOO0ooiiLliio );
 OoOOIil0oLiOILOIIIlIli000O0il000I <= OO0o0l0ioiI0oo0oiOL00LooiIIoli00o;
 end
 else begin
 OiILLloIOIIolIio00l00OLOLLIlLoO0o <= 1'b0;
 OLl0l0oIIoi00000IiiloiLi0OoloLi0L <= 3'b0;
 OL0Ioll0l0OiIOliOLollLOil000o0iol <= 1'b0;
 OoOOIil0oLiOILOIIIlIli000O0il000I <= 64'b0;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(Olo0I0OOli0Oii0IoOOLloiiliollIolO == SEARCH) begin
 if(OLOIl0loioiIllIlOlOLiOO0ooiiLliio & OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL) OLi00LI00i0LIIiO0olIo00Liii0ILLii <= 1'b1;
 end
 else OLi00LI00i0LIIiO0olIo00Liii0ILLii <= 5'b0;
 wire OiIIloOooI0IoLLO0ILlIi0LoiiLl00OO;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo <= 1'b0;
 else if((Olo0I0OOli0Oii0IoOOLloiiliollIolO == PAYLOAD_OUT) && O0L00liiLLLiiL00OlOoOilOOiil00LIl) O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo <= 1'b1;
 else if((Olo0I0OOli0Oii0IoOOLloiiliollIolO == SEARCH) && OLOIl0loioiIllIlOlOLiOO0ooiiLliio) O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo <= 1'b1;
 assign OiIIloOooI0IoLLO0ILlIi0LoiiLl00OO = O0iliOIiiLOoi0OiOOoiooIOiilL0OoIo || ((Olo0I0OOli0Oii0IoOOLloiiliollIolO == PAYLOAD_OUT) && O0L00liiLLLiiL00OlOoOilOOiil00LIl) || ((Olo0I0OOli0Oii0IoOOLloiiliollIolO == SEARCH) && OLOIl0loioiIllIlOlOLiOO0ooiiLliio);
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) begin
 O0LIllilOiLIoilOlLiOio0LiILlllLiI <= OoIlOoIlIooO0lIIooIoillLl0O0OLlol ;
 OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO <= OOLOOIi000oLlOiO0LLiIIIoIIO0ILool;
 end
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) OoiillIIi0O00lLlIOOiO0OOii0LiLiLO <= 'd0;
 else if(OlOiLILOlooo00OLIILLiOioIlO0lLi0l) OoiillIIi0O00lLlIOOiO0OOii0LiLiLO <= OoiillIIi0O00lLlIOOiO0OOii0LiLiLO + 1'b1;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) O0li0Illi0oOollo0ooOoIiolOoio0iiL <= 64'd0;
 else if(OiILLloIOIIolIio00l00OLOLLIlLoO0o&&OL0Ioll0l0OiIOliOLollLOil000o0iol) O0li0Illi0oOollo0ooOoIiolOoio0iiL <= O0li0Illi0oOollo0ooOoIiolOoio0iiL + 1'b1;
 always @(posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(!OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI) OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil <= 32'd0;
 else if(OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL &&(OillLLIloOooLolooI0oiLLOO0LOoliio == 8'd2)&&(OO0o0l0ioiI0oo0oiOL00LooiIIoli00o[7:0]==8'h06)) OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil <= OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil + 1'b1;
 endmodule
 module OOLIoOio0I0i0lliO0OoolLLLLIoLLLlI ( O0oLi000Lo0oO0oLLoIOllIlo0iOoILio, OiloLLIoolOIiOiOoo00L0I0IOio0lI0L, Ol00oIollLiioLLLoiOiolOL00iiOlIoo, OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI, OOLOlOo0000iOi0OLOolloLo0iL0iooIi, OL0IIIOOo0000OLoOiO00iiO0lLolLIoO, OIoII0liiOiiO0Lo0illI0iOOI0ll000I, OlOiLILOlooo00OLIILLiOioIlO0lLi0l, OiiillOL0OL0oI0O0liIlLIIOL0iLLIli, OlOlLl00OLLOO0ooloIoIli0IIoOLIlOo, OOlOiil0loi0LllL0oOLI00OLoil0l0Ii, OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl, Olli0loIii0llI00IoOlO0iloLI0oOLOI, OloOoiioIil00OoLilIliO00IiiillI0I, O00iLoILoLlOOOolIiiiIOOIlILliLIO0, OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl, OlLILLOo0IOoilLOO0OlLiioiiioi0IlL, OL0Ioll0l0OiIOliOLollLOil000o0iol, OoOOIil0oLiOILOIIIlIli000O0il000I, OiILLloIOIIolIio00l00OLOLLIlLoO0o, OLl0l0oIIoi00000IiiloiLi0OoloLi0L, O0LIllilOiLIoilOlLiOio0LiILlllLiI, OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO, OiIoiiOIOOi0OLILo0oIOOioO0IioLI00, OLll00OOliOil0O0iLlIooLOLooIIlI0o, OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0, OOLIiil0IlIllLollIl0LIilliOI0iolo, OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 , OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI , OolIOLOooiLLIllI0LOLIolllLoilolIl , O0IOooLliOlIllOliILoolIIoIiO0Ilol , OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI , OilOOo00lLiOOoiO0ii0oo0oOliOollii , OLo0oiiL0ooIliO0I0illLoILiiIoIoOI , OO0liOO0iOOIioool0OoLliiiI0l0ilOo , OiIOLi00lOILlOOL0oLLloL0io0LoIoOL , OIloLiiOL00oilLo0iiILoOOll0lIlIlO, OoiillIIi0O00lLlIOOiO0OOii0LiLiLO, OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil, O0li0Illi0oOollo0ooOoIiolOoio0iiL );
 input O0oLi000Lo0oO0oLLoIOllIlo0iOoILio;
 input OiloLLIoolOIiOiOoo00L0I0IOio0lI0L;
 input Ol00oIollLiioLLLoiOiolOL00iiOlIoo;
 input OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI;
 input OOLOlOo0000iOi0OLOolloLo0iL0iooIi;
 input OL0IIIOOo0000OLoOiO00iiO0lLolLIoO;
 input [31:0] OIoII0liiOiiO0Lo0illI0iOOI0ll000I;
 input OlOiLILOlooo00OLIILLiOioIlO0lLi0l;
 input OiiillOL0OL0oI0O0liIlLIIOL0iLLIli;
 input [1:0] OlOlLl00OLLOO0ooloIoIli0IIoOLIlOo;
 input [31:0] OOlOiil0loi0LllL0oOLI00OLoil0l0Ii;
 input [31:0] OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl;
 output [15:0] Olli0loIii0llI00IoOlO0iloLI0oOLOI;
 output [15:0] OloOoiioIil00OoLilIliO00IiiillI0I;
 output [31:0] O00iLoILoLlOOOolIiiiIOOIlILliLIO0;
 output [31:0] OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl;
 input OlLILLOo0IOoilLOO0OlLiioiiioi0IlL;
 output OL0Ioll0l0OiIOliOLollLOil000o0iol;
 output [63:0] OoOOIil0oLiOILOIIIlIli000O0il000I;
 output OiILLloIOIIolIio00l00OLOLLIlLoO0o;
 output [3:0] OLl0l0oIIoi00000IiiloiLi0OoloLi0L;
 output O0LIllilOiLIoilOlLiOio0LiILlllLiI;
 output [2:0] OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO;
 output [15:0] OiIoiiOIOOi0OLILo0oIOOioO0IioLI00;
 input [31:0] OLll00OOliOil0O0iLlIooLOLooIIlI0o;
 input [31:0] OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0;
 input [4:0] OOLIiil0IlIllLollIl0LIilliOI0iolo;
 input OLOILlOloOoi0OO0oLOOlo0iiIoioilL0 ;
 input [3:0] OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI ;
 input [15:0] OolIOLOooiLLIllI0LOLIolllLoilolIl ;
 input [ 5:0] O0IOooLliOlIllOliILoolIIoIiO0Ilol ;
 input [5:0] OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI ;
 input OilOOo00lLiOOoiO0ii0oo0oOliOollii ;
 input [31:0 ] OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ;
 input [31:0 ] OO0liOO0iOOIioool0OoLliiiI0l0ilOo ;
 input OiIOLi00lOILlOOL0oLLloL0io0LoIoOL ;
 input [31:0] OIloLiiOL00oilLo0iiILoOOll0lIlIlO;
 output [63:0] OoiillIIi0O00lLlIOOiO0OOii0LiLiLO;
 output [31:0] OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil;
 output [63:0] O0li0Illi0oOollo0ooOoIiolOoio0iiL;
 wire OiLOOl0Lo0OI0loiloLIoLLiIoLILliLi;
 wire [63:0] OLLOooI0ILL00ILloiliILLLiioooLliI;
 wire OiLOiiLLloIliLlOLI00O0iiioooLloIO;
 wire Oool000Ii0llLOoILOIloiO0oIlIoL0oO;
 wire [2:0] OLIo0lIO0IL0LlO0LIOoolOIlI0OOl0iL;
 wire OOii0olOiiL0loIO0oiliLOIiOOL0Lol0;
 wire OoLOOii0LIioLOolIiLLOIIOiiIOLlool;
 reg [11:0] O0ILlL0loOoLO0ooILIoOoiIILooIooOo;
 reg [11:0] OLIIli0LOiLIILloiolioLilOoOL00iOI;
 always @ (posedge Ol00oIollLiioLLLoiOiolOL00iiOlIoo) if(OOLOlOo0000iOi0OLOolloLo0iL0iooIi) O0ILlL0loOoLO0ooILIoOoiIILooIooOo <= 12'h0;
 else O0ILlL0loOoLO0ooILIoOoiIILooIooOo <= {O0ILlL0loOoLO0ooILIoOoiIILooIooOo[10:0],1'b1};
 assign OoLOOii0LIioLOolIiLLOIIOiiIOLlool = O0ILlL0loOoLO0ooILIoOoiIILooIooOo[11];
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) if(OOLOlOo0000iOi0OLOolloLo0iL0iooIi) OLIIli0LOiLIILloiolioLilOoOL00iOI <= 12'h0;
 else OLIIli0LOiLIILloiolioLilOoOL00iOI <= {OLIIli0LOiLIILloiolioLilOoOL00iOI[10:0],1'b1};
 assign OOii0olOiiL0loIO0oiliLOIiOOL0Lol0 = OLIIli0LOiLIILloiolioLilOoOL00iOI[11];
 OO0iLlLLlL0LII000oOLLILOliLLO00iL u_wrapper_mac_rx_fifo ( .O0oLi000Lo0oO0oLLoIOllIlo0iOoILio (O0oLi000Lo0oO0oLLoIOllIlo0iOoILio), .OiloLLIoolOIiOiOoo00L0I0IOio0lI0L (OiloLLIoolOIiOiOoo00L0I0IOio0lI0L&&OOii0olOiiL0loIO0oiliLOIiOOL0Lol0), .OIoII0liiOiiO0Lo0illI0iOOI0ll000I (OIoII0liiOiiO0Lo0illI0iOOI0ll000I), .OoIO00ILLOLIoiI00IoOiIioILOLO0iOO (OlOlLl00OLLOO0ooloIoIli0IIoOLIlOo), .OL0IIIOOo0000OLoOiO00iiO0lLolLIoO (OL0IIIOOo0000OLoOiO00iiO0lLolLIoO), .OlOiLILOlooo00OLIILLiOioIlO0lLi0l (OlOiLILOlooo00OLIILLiOioIlO0lLi0l), .OiiillOL0OL0oI0O0liIlLIIOL0iLLIli (OiiillOL0OL0oI0O0liIlLIIOL0iLLIli), .OOIoloilOiLOIOliIOI0oli0oiiiILlI0 (Ol00oIollLiioLLLoiOiolOL00iiOlIoo), .OlLILLOo0IOoilLOO0OlLiioiiioi0IlL (OlLILLOo0IOoilLOO0OlLiioiiioi0IlL), .OIOoIILIooOiOOLIOIll0IIl0LolIiilo (OLLOooI0ILL00ILloiliILLLiioooLliI), .OIliIOoLL0OI0l0i0iiiOLi0lLLilLiOI (OLIo0lIO0IL0LlO0LIOoolOIlI0OOl0iL), .OiLIIiiIooi0LllOiIilO0LIi0l00i0iL (OiLOOl0Lo0OI0loiloLIoLLiIoLILliLi), .O0OlLLoiol0OLiii0LO0oolloLLoolIli (OiLOiiLLloIliLlOLI00O0iiioooLloIO), .Oi0iOLLIoO00iLLLoOOOo0LIoLlII00II (Oool000Ii0llLOoILOIloiO0oIlIoL0oO) );
 OoILi0OOLIloI0O0lO0lOLo0iLlO0o0oo OiLooiOOioILOo0lLlli0Liol0iOo00ol( .Ol00oIollLiioLLLoiOiolOL00iiOlIoo (Ol00oIollLiioLLLoiOiolOL00iiOlIoo), .OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI (OloIiOlOoILlLoLOiLIIIIoloOoIiLoiI&&OoLOOii0LIioLOolIiLLOIIOiiIOLlool), .OiLIiLoILI0LiLOlLIoOolOolIIlOIllI (OOLIiil0IlIllLollIl0LIilliOI0iolo), .OiiiIllliL0oLoOIliliIilLiollooiII( OLOILlOloOoi0OO0oLOOlo0iiIoioilL0) , .OI0ioooOlLlIoLiL0IO0oOII0OlLiOo0I (OloO0OIiOLi0LlIlILiOoO0iiLooo0LiI), .O0lOOlIOlIo0IILillLi0liOLlO00OILL (OolIOLOooiLLIllI0LOLIolllLoilolIl), .OILLO0olLiLlOoOolOloOOLiliIIiIOLO (O0IOooLliOlIllOliILoolIIoIiO0Ilol), .OIiOoioOIOoLIOO0OLioll0I0IIiIoOOi (OOL0o0IoOoIooIL0Ool0l0iOIIlIliOlI), .OOIOlI0OolOlLlOOIii0ioo00iio0IIil (OilOOo00lLiOOoiO0ii0oo0oOliOollii), .OIloLiiOL00oilLo0iiILoOOll0lIlIlO (OIloLiiOL00oilLo0iiILoOOll0lIlIlO), .OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ( OLo0oiiL0ooIliO0I0illLoILiiIoIoOI ), .OO0liOO0iOOIioool0OoLliiiI0l0ilOo (OO0liOO0iOOIioool0OoLliiiI0l0ilOo ), .OiIOLi00lOILlOOL0oLLloL0io0LoIoOL (OiIOLi00lOILlOOL0oLLloL0io0LoIoOL), .OoLIIO0Oi0oOO0o0LOLiLIlLlLloIoIiL (OiLOOl0Lo0OI0loiloLIoLLiIoLILliLi), .OO0o0l0ioiI0oo0oiOL00LooiIIoli00o (OLLOooI0ILL00ILloiliILLLiioooLliI), .OollLiiii0o0lIiIiL0OL0OLiLllLL0I0 (OiLOiiLLloIliLlOLI00O0iiioooLloIO), .OoIlOoIlIooO0lIIooIoillLl0O0OLlol (Oool000Ii0llLOoILOIloiO0oIlIoL0oO), .OOLOOIi000oLlOiO0LLiIIIoIIO0ILool (OLIo0lIO0IL0LlO0LIOoolOIlI0OOl0iL), .OOlOiil0loi0LllL0oOLI00OLoil0l0Ii (OOlOiil0loi0LllL0oOLI00OLoil0l0Ii), .OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl (OLoLOOIlolLI0iOLiIlLol0lLLoolOiLl), .Olli0loIii0llI00IoOlO0iloLI0oOLOI (Olli0loIii0llI00IoOlO0iloLI0oOLOI), .OloOoiioIil00OoLilIliO00IiiillI0I (OloOoiioIil00OoLilIliO00IiiillI0I), .O00iLoILoLlOOOolIiiiIOOIlILliLIO0 (O00iLoILoLlOOOolIiiiIOOIlILliLIO0), .OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl (OLO00Ooiio0IoiLiOLIoIOIiOi0IooiOl), .OL0Ioll0l0OiIOliOLollLOil000o0iol (OL0Ioll0l0OiIOliOLollLOil000o0iol), .OoOOIil0oLiOILOIIIlIli000O0il000I (OoOOIil0oLiOILOIIIlIli000O0il000I), .OiILLloIOIIolIio00l00OLOLLIlLoO0o (OiILLloIOIIolIio00l00OLOLLIlLoO0o), .OLl0l0oIIoi00000IiiloiLi0OoloLi0L (OLl0l0oIIoi00000IiiloiLi0OoloLi0L), .O0LIllilOiLIoilOlLiOio0LiILlllLiI (O0LIllilOiLIoilOlLiOio0LiILlllLiI), .OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO (OiOOLLIllIOoILiIOlLLLIiLlI0OIOLoO), .OiIoiiOIOOi0OLILo0oIOOioO0IioLI00 (OiIoiiOIOOi0OLILo0oIOOioO0IioLI00), .OoiillIIi0O00lLlIOOiO0OOii0LiLiLO (OoiillIIi0O00lLlIOOiO0OOii0LiLiLO), .OLll00OOliOil0O0iLlIooLOLooIIlI0o (OLll00OOliOil0O0iLlIooLOLooIIlI0o), .OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0(OoOl0LLiiLiiLIO00O0O0ioLo0OIiioI0), .OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil (OOIILlLoiiLOoI0iOiLLoL0ilIOiLlLil), .O0li0Illi0oOollo0ooOoIiolOoio0iiL (O0li0Illi0oOollo0ooOoIiolOoio0iiL) );
 endmodule
 module OO0iLlLLlL0LII000oOLLILOliLLO00iL( O0oLi000Lo0oO0oLLoIOllIlo0iOoILio, OiloLLIoolOIiOiOoo00L0I0IOio0lI0L, OIoII0liiOiiO0Lo0illI0iOOI0ll000I, OoIO00ILLOLIoiI00IoOiIioILOLO0iOO, OL0IIIOOo0000OLoOiO00iiO0lLolLIoO, OlOiLILOlooo00OLIILLiOioIlO0lLi0l, OiiillOL0OL0oI0O0liIlLIIOL0iLLIli, OOIoloilOiLOIOliIOI0oli0oiiiILlI0, OlLILLOo0IOoilLOO0OlLiioiiioi0IlL, OIOoIILIooOiOOLIOIll0IIl0LolIiilo, OIliIOoLL0OI0l0i0iiiOLi0lLLilLiOI, OiLIIiiIooi0LllOiIilO0LIi0l00i0iL, O0OlLLoiol0OLiii0LO0oolloLLoolIli, Oi0iOLLIoO00iLLLoOOOo0LIoLlII00II );
 input O0oLi000Lo0oO0oLLoIOllIlo0iOoILio;
 input OiloLLIoolOIiOiOoo00L0I0IOio0lI0L;
 input [31:0] OIoII0liiOiiO0Lo0illI0iOOI0ll000I;
 input [1:0] OoIO00ILLOLIoiI00IoOiIioILOLO0iOO;
 input OL0IIIOOo0000OLoOiO00iiO0lLolLIoO;
 input OlOiLILOlooo00OLIILLiOioIlO0lLi0l;
 input OiiillOL0OL0oI0O0liIlLIIOL0iLLIli;
 input OOIoloilOiLOIOliIOI0oli0oiiiILlI0;
 input OlLILLOo0IOoilLOO0OlLiioiiioi0IlL;
 output [63:0] OIOoIILIooOiOOLIOIll0IIl0LolIiilo;
 output [2:0] OIliIOoLL0OI0l0i0iiiOLi0lLLilLiOI;
 output OiLIIiiIooi0LllOiIilO0LIi0l00i0iL;
 output O0OlLLoiol0OLiii0LO0oolloLLoolIli;
 output Oi0iOLLIoO00iLLLoOOOo0LIoLlII00II;
 wire OoLoiIlIlOLo0IiO0lOolLLoo0I0Io0IO;
 wire OIOlO0iOoIL0OoO0oIoilooILI00iIIOL;
 wire [69:0] OloLIlO0L00loIO0ol0ioIIoooLioiLlo;
 wire [69:0] OIiiIlI0oIOIIolIoLoLliOoLlIloIioi;
 reg OlOo0OO0lo0ooOoII0llOlOIoOLoIoilo;
 wire OlilL0OLLI0l0LOLOLOl0iLolIolOLLoI;
 reg O0l0liI00iI0ooi0o0OL00oo0o0iIILlO;
 reg [35:0] Oil0OLI0o0l0iIlL0oooIIOoO00LoLIiI;
 reg [2:0] O0LIIIILLiOOlOOOlLoo0iOoLio0iO0Il;
 reg [63:0] OIlIOoI0oliLooOIIOOLLolooloL0LiLl;
 wire [1:0] O00iLLLLlOl00oI0loO0OllooooiILolo;
 reg OoloIOILLOlLIOIolIi0iIllLi0ilioLL;
 reg O0LlO00lILOIOlil0IILLlIiooio0iILO;
 assign O00iLLLLlOl00oI0loO0OllooooiILolo = 3'd4 - OoIO00ILLOLIoiI00IoOiIioILOLO0iOO;
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) if(!OiloLLIoolOIiOiOoo00L0I0IOio0lI0L) O0l0liI00iI0ooi0o0OL00oo0o0iIILlO <= 1'b0;
 else if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO & OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) O0l0liI00iI0ooi0o0OL00oo0o0iIILlO <= 1'b0;
 else if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO) O0l0liI00iI0ooi0o0OL00oo0o0iIILlO <= ~O0l0liI00iI0ooi0o0OL00oo0o0iIILlO;
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO && !O0l0liI00iI0ooi0o0OL00oo0o0iIILlO) Oil0OLI0o0l0iIlL0oooIIOoO00LoLIiI <= {OlOiLILOlooo00OLIILLiOioIlO0lLi0l,OiiillOL0OL0oI0O0liIlLIIOL0iLLIli,O00iLLLLlOl00oI0loO0OllooooiILolo,OIoII0liiOiiO0Lo0illI0iOOI0ll000I};
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO && OiiillOL0OL0oI0O0liIlLIIOL0iLLIli && O0l0liI00iI0ooi0o0OL00oo0o0iIILlO) O0LIIIILLiOOlOOOlLoo0iOoLio0iO0Il <= {1'b0,O00iLLLLlOl00oI0loO0OllooooiILolo};
 else if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO && OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) O0LIIIILLiOOlOOOlLoo0iOoLio0iO0Il <= {1'b1,O00iLLLLlOl00oI0loO0OllooooiILolo};
 else O0LIIIILLiOOlOOOlLoo0iOoLio0iO0Il <= 3'b0;
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO && OiiillOL0OL0oI0O0liIlLIIOL0iLLIli && O0l0liI00iI0ooi0o0OL00oo0o0iIILlO) OIlIOoI0oliLooOIIOOLLolooloL0LiLl <= {Oil0OLI0o0l0iIlL0oooIIOoO00LoLIiI[31:0],OIoII0liiOiiO0Lo0illI0iOOI0ll000I};
 else if(OL0IIIOOo0000OLoOiO00iiO0lLolLIoO && OiiillOL0OL0oI0O0liIlLIIOL0iLLIli) OIlIOoI0oliLooOIIOOLLolooloL0LiLl <= {OIoII0liiOiiO0Lo0illI0iOOI0ll000I,32'b0};
 else OIlIOoI0oliLooOIIOOLLolooloL0LiLl <= {Oil0OLI0o0l0iIlL0oooIIOoO00LoLIiI[31:0],OIoII0liiOiiO0Lo0illI0iOOI0ll000I};
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) begin
 if(!OiloLLIoolOIiOiOoo00L0I0IOio0lI0L) OlOo0OO0lo0ooOoII0llOlOIoOLoIoilo <= 1'b0;
 else OlOo0OO0lo0ooOoII0llOlOIoOLoIoilo <= OL0IIIOOo0000OLoOiO00iiO0lLolLIoO & O0l0liI00iI0ooi0o0OL00oo0o0iIILlO | OL0IIIOOo0000OLoOiO00iiO0lLolLIoO & OiiillOL0OL0oI0O0liIlLIIOL0iLLIli;
 end
 always @ (posedge O0oLi000Lo0oO0oLLoIOllIlo0iOoILio) if(!OiloLLIoolOIiOiOoo00L0I0IOio0lI0L) begin
 O0LlO00lILOIOlil0IILLlIiooio0iILO <= 1'b0;
 OoloIOILLOlLIOIolIi0iIllLi0ilioLL <= 1'b0;
 end
 else begin
 O0LlO00lILOIOlil0IILLlIiooio0iILO <= Oil0OLI0o0l0iIlL0oooIIOoO00LoLIiI[35];
 OoloIOILLOlLIOIolIi0iIllLi0ilioLL <= OiiillOL0OL0oI0O0liIlLIIOL0iLLIli;
 end
 assign OloLIlO0L00loIO0ol0ioIIoooLioiLlo = {1'b0,O0LlO00lILOIOlil0IILLlIiooio0iILO,OoloIOILLOlLIOIolIi0iIllLi0ilioLL,O0LIIIILLiOOlOOOlLoo0iOoLio0iO0Il,OIlIOoI0oliLooOIIOOLLolooloL0LiLl};
 assign OlilL0OLLI0l0LOLOLOl0iLolIolOLLoI = !OIOlO0iOoIL0OoO0oIoilooILI00iIIOL && OlLILLOo0IOoilLOO0OlLiioiiioi0IlL;
 assign OIOoIILIooOiOOLIOIll0IIl0LolIiilo = OIiiIlI0oIOIIolIoLoLliOoLlIloIioi[63:0];
 assign OIliIOoLL0OI0l0i0iiiOLi0lLLilLiOI = OIiiIlI0oIOIIolIoLoLliOoLlIloIioi[66:64];
 assign O0OlLLoiol0OLiii0LO0oolloLLoolIli = OIiiIlI0oIOIIolIoLoLliOoLlIloIioi[68];
 assign Oi0iOLLIoO00iLLLoOOOo0LIoLlII00II = OIiiIlI0oIOIIolIoLoLliOoLlIloIioi[67];
 assign OiLIIiiIooi0LllOiIilO0LIi0l00i0iL = OlilL0OLLI0l0LOLOLOl0iLolIolOLLoI;
 mac_rx_fifo OO0iLlLLlL0LII000oOLLILOliLLO00iL( .data (OloLIlO0L00loIO0ol0ioIIoooLioiLlo), .wrreq (OlOo0OO0lo0ooOoII0llOlOIoOLoIoilo), .rdreq (OlilL0OLLI0l0LOLOLOl0iLolIolOLLoI), .wrclk (O0oLi000Lo0oO0oLLoIOllIlo0iOoILio), .rdclk (OOIoloilOiLOIOliIOI0oli0oiiiILlI0), .q (OIiiIlI0oIOIIolIoLoLliOoLlIloIioi), .rdempty (OIOlO0iOoIL0OoO0oIoilooILI00iIIOL), .wrfull (OoLoiIlIlOLo0IiO0lOolLLoo0I0Io0IO) );
 endmodule
 